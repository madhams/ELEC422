magic
tech scmos
timestamp 1681772484
<< nwell >>
rect -1 3654 41 3695
rect 285 3652 330 3692
rect 599 3654 645 3693
rect 914 3651 953 3687
rect 1202 3661 1243 3695
rect 1516 3658 1550 3691
rect 1804 3658 1846 3698
rect 2100 3642 2139 3681
rect 2404 3644 2450 3692
rect 2692 3641 2737 3686
rect -1017 2631 -982 2669
rect 3727 2625 3753 2657
rect -1015 2337 -978 2372
rect 3725 2342 3760 2374
rect -1020 2027 -989 2060
rect 3719 2030 3748 2063
rect -1015 1735 -982 1769
rect 3730 1742 3760 1770
rect -1018 1445 -986 1478
rect 3736 1432 3764 1459
rect -1030 1125 -1000 1157
rect 3723 1142 3756 1174
rect -1016 830 -989 854
rect 3728 849 3750 870
rect -1020 538 -996 563
rect 3731 545 3756 570
rect -1023 245 -998 269
rect 3726 240 3752 268
rect -1024 -67 -993 -38
rect 3728 -65 3756 -35
rect 14 -1069 40 -1044
rect 311 -1078 343 -1050
rect 609 -1079 639 -1052
rect 914 -1072 941 -1046
rect 1205 -1055 1224 -1038
rect 1511 -1076 1536 -1053
rect 1816 -1074 1846 -1048
rect 2110 -1091 2138 -1067
rect 2418 -1094 2446 -1066
rect 2713 -1085 2736 -1061
<< polysilicon >>
rect 3598 3774 3853 3775
rect -1108 3482 -132 3750
rect 2910 3514 3853 3774
rect -1108 2818 -828 3482
rect 3598 2836 3853 3514
rect -70 2644 2833 2761
rect -68 -156 1185 -16
rect 1249 -150 2750 -10
rect -1095 -917 -816 -222
rect 3570 -917 3853 -278
rect -1096 -1186 -164 -917
rect 2890 -1180 3853 -917
rect 2890 -1191 3851 -1180
<< metal1 >>
rect 3598 3774 3853 3775
rect -1108 3482 -132 3750
rect 2910 3514 3853 3774
rect -1108 2818 -828 3482
rect 3598 2836 3853 3514
rect 1523 2775 1527 2789
rect -97 2771 199 2775
rect 203 2771 499 2775
rect 503 2771 799 2775
rect 803 2771 1347 2775
rect 1351 2771 1699 2775
rect 1703 2771 1999 2775
rect 2003 2771 2299 2775
rect 2303 2771 2599 2775
rect 2603 2771 2844 2775
rect -101 2476 -97 2771
rect -70 2644 2833 2761
rect 14 2607 2722 2627
rect 38 2583 2698 2603
rect 38 2567 2698 2573
rect 666 2526 669 2535
rect 682 2533 692 2536
rect 1162 2533 1172 2536
rect 1492 2533 1500 2536
rect 1604 2533 1612 2536
rect 1660 2533 1668 2536
rect 1722 2533 1780 2536
rect 1796 2533 1805 2536
rect 1826 2526 1829 2545
rect 1906 2543 1916 2546
rect 1964 2543 1973 2546
rect 1970 2536 1973 2543
rect 1836 2533 1853 2536
rect 1924 2533 1941 2536
rect 1970 2533 1988 2536
rect 2034 2533 2044 2536
rect 2098 2533 2116 2536
rect 204 2523 229 2526
rect 300 2523 317 2526
rect 604 2523 629 2526
rect 660 2523 669 2526
rect 676 2523 693 2526
rect 708 2523 725 2526
rect 812 2523 828 2526
rect 1012 2523 1037 2526
rect 1068 2523 1077 2526
rect 1084 2523 1100 2526
rect 1114 2523 1132 2526
rect 1156 2523 1173 2526
rect 1194 2523 1204 2526
rect 1316 2523 1333 2526
rect 1524 2523 1533 2526
rect 1698 2523 1772 2526
rect 1804 2523 1813 2526
rect 1820 2523 1829 2526
rect 690 2515 693 2523
rect 1114 2515 1117 2523
rect 1850 2506 1853 2533
rect 1890 2523 1900 2526
rect 1938 2525 1941 2533
rect 2186 2526 2189 2535
rect 2236 2533 2253 2536
rect 2266 2526 2269 2535
rect 2314 2533 2324 2536
rect 2378 2533 2388 2536
rect 1964 2523 1973 2526
rect 2004 2523 2028 2526
rect 2034 2523 2060 2526
rect 2180 2523 2189 2526
rect 2220 2523 2269 2526
rect 2290 2523 2308 2526
rect 2396 2523 2405 2526
rect 2420 2523 2428 2526
rect 2460 2523 2476 2526
rect 2490 2525 2493 2536
rect 2564 2533 2629 2536
rect 2538 2523 2548 2526
rect 1978 2513 1988 2516
rect 2292 2513 2301 2516
rect 2316 2513 2325 2516
rect 1850 2503 1876 2506
rect 2844 2476 2848 2771
rect -101 2176 -97 2472
rect 14 2467 2722 2473
rect 714 2433 724 2436
rect 1762 2433 1804 2436
rect 1938 2433 1948 2436
rect 2546 2433 2556 2436
rect 676 2423 685 2426
rect 882 2423 892 2426
rect 1034 2416 1037 2425
rect 1186 2416 1189 2425
rect 1778 2423 1788 2426
rect 1844 2423 1869 2426
rect 2018 2423 2028 2426
rect 2042 2423 2052 2426
rect 2364 2423 2373 2426
rect 2530 2423 2540 2426
rect 2570 2423 2580 2426
rect 124 2413 149 2416
rect 180 2413 189 2416
rect 196 2413 205 2416
rect 244 2413 261 2416
rect 66 2403 76 2406
rect 202 2405 205 2413
rect 258 2405 261 2413
rect 330 2413 340 2416
rect 346 2413 357 2416
rect 402 2413 412 2416
rect 474 2413 484 2416
rect 522 2413 532 2416
rect 538 2413 565 2416
rect 636 2413 645 2416
rect 674 2413 692 2416
rect 330 2405 333 2413
rect 346 2405 349 2413
rect 354 2403 372 2406
rect 402 2405 405 2413
rect 420 2403 437 2406
rect 522 2405 525 2413
rect 538 2406 541 2413
rect 538 2405 549 2406
rect 540 2403 549 2405
rect 634 2403 652 2406
rect 714 2403 717 2414
rect 762 2413 772 2416
rect 786 2405 789 2416
rect 834 2413 844 2416
rect 868 2413 885 2416
rect 948 2413 973 2416
rect 1010 2413 1020 2416
rect 1034 2413 1052 2416
rect 1100 2413 1125 2416
rect 1156 2413 1165 2416
rect 1186 2413 1204 2416
rect 1274 2413 1300 2416
rect 1314 2413 1332 2416
rect 1426 2413 1452 2416
rect 1490 2413 1508 2416
rect 1546 2413 1572 2416
rect 1722 2413 1740 2416
rect 1818 2413 1828 2416
rect 1850 2413 1884 2416
rect 842 2403 852 2406
rect 1218 2403 1228 2406
rect 1276 2403 1285 2406
rect 1418 2403 1428 2406
rect 1482 2403 1492 2406
rect 1602 2403 1620 2406
rect 1730 2403 1748 2406
rect 1844 2403 1861 2406
rect 1906 2403 1925 2406
rect 1938 2403 1941 2414
rect 1980 2413 2029 2416
rect 2036 2413 2053 2416
rect 2074 2413 2092 2416
rect 2098 2413 2108 2416
rect 2186 2413 2212 2416
rect 2074 2405 2077 2413
rect 2274 2406 2277 2414
rect 2324 2413 2341 2416
rect 2412 2413 2436 2416
rect 2460 2413 2477 2416
rect 2260 2403 2277 2406
rect 2338 2405 2341 2413
rect 2498 2406 2501 2414
rect 2524 2413 2533 2416
rect 2364 2403 2373 2406
rect 2434 2403 2444 2406
rect 2466 2403 2501 2406
rect 2626 2403 2636 2406
rect 1890 2393 1908 2396
rect 2300 2393 2309 2396
rect 38 2367 2698 2373
rect 642 2343 652 2346
rect 1474 2343 1493 2346
rect 1866 2343 1876 2346
rect 2018 2336 2021 2345
rect 66 2333 76 2336
rect 186 2326 189 2335
rect 202 2326 205 2335
rect 242 2333 268 2336
rect 282 2326 285 2335
rect 490 2326 493 2335
rect 636 2333 645 2336
rect 660 2333 677 2336
rect 698 2333 724 2336
rect 124 2323 149 2326
rect 180 2323 189 2326
rect 196 2323 205 2326
rect 276 2323 285 2326
rect 292 2323 317 2326
rect 490 2323 500 2326
rect 610 2323 628 2326
rect 674 2325 677 2333
rect 706 2323 732 2326
rect 738 2325 741 2336
rect 748 2333 757 2336
rect 770 2325 773 2336
rect 794 2333 804 2336
rect 828 2333 861 2336
rect 940 2333 973 2336
rect 1092 2333 1141 2336
rect 1162 2333 1276 2336
rect 1300 2333 1317 2336
rect 1468 2333 1508 2336
rect 1556 2333 1565 2336
rect 1572 2333 1581 2336
rect 1642 2333 1668 2336
rect 1716 2333 1725 2336
rect 834 2313 868 2316
rect 874 2306 877 2325
rect 970 2323 973 2333
rect 1042 2323 1084 2326
rect 1562 2325 1565 2333
rect 1658 2323 1676 2326
rect 1682 2323 1700 2326
rect 1738 2325 1741 2336
rect 1770 2333 1780 2336
rect 1796 2333 1805 2336
rect 1826 2333 1844 2336
rect 1884 2333 1909 2336
rect 2012 2333 2021 2336
rect 2050 2333 2068 2336
rect 2202 2333 2212 2336
rect 2242 2333 2252 2336
rect 2258 2333 2316 2336
rect 1762 2323 1772 2326
rect 1804 2323 1813 2326
rect 1898 2323 1908 2326
rect 1956 2324 1980 2327
rect 2044 2323 2053 2326
rect 2076 2323 2085 2326
rect 2204 2323 2213 2326
rect 2260 2323 2277 2326
rect 2330 2325 2333 2336
rect 2340 2333 2357 2336
rect 2370 2325 2373 2336
rect 2466 2333 2476 2336
rect 2586 2333 2596 2336
rect 2644 2333 2653 2336
rect 1058 2313 1076 2316
rect 1300 2313 1309 2316
rect 1954 2313 1964 2316
rect 2082 2313 2092 2316
rect 2116 2313 2125 2316
rect 2388 2313 2405 2316
rect 2402 2306 2405 2313
rect 2418 2306 2421 2325
rect 2450 2323 2484 2326
rect 2548 2324 2564 2327
rect 2620 2323 2669 2326
rect 2436 2313 2469 2316
rect 770 2303 780 2306
rect 850 2303 877 2306
rect 1948 2303 1965 2306
rect 2362 2303 2380 2306
rect 2402 2303 2421 2306
rect 2562 2303 2572 2306
rect 14 2267 2722 2273
rect 842 2233 876 2236
rect 1476 2233 1501 2236
rect 1858 2233 1876 2236
rect 2458 2233 2468 2236
rect 2498 2233 2516 2236
rect 842 2223 860 2226
rect 884 2223 933 2226
rect 1298 2216 1301 2225
rect 1458 2223 1468 2226
rect 1538 2216 1541 2225
rect 1692 2223 1717 2226
rect 1842 2223 1860 2226
rect 2250 2216 2253 2225
rect 2506 2217 2509 2226
rect 74 2213 84 2216
rect 100 2213 109 2216
rect 276 2213 285 2216
rect 292 2213 317 2216
rect 322 2213 332 2216
rect 66 2203 76 2206
rect 258 2203 268 2206
rect 338 2205 341 2216
rect 428 2213 437 2216
rect 346 2203 356 2206
rect 388 2203 413 2206
rect 434 2205 437 2213
rect 450 2203 460 2206
rect 490 2203 508 2206
rect 540 2203 581 2206
rect 586 2205 589 2216
rect 596 2213 613 2216
rect 652 2213 661 2216
rect 674 2213 708 2216
rect 820 2213 829 2216
rect 836 2213 853 2216
rect 996 2213 1013 2216
rect 1018 2213 1028 2216
rect 1210 2213 1236 2216
rect 1298 2213 1316 2216
rect 1516 2213 1541 2216
rect 1620 2213 1653 2216
rect 1684 2213 1717 2216
rect 1756 2213 1765 2216
rect 1770 2213 1780 2216
rect 1812 2213 1820 2216
rect 610 2206 613 2213
rect 610 2203 628 2206
rect 658 2205 661 2213
rect 682 2203 700 2206
rect 724 2203 773 2206
rect 780 2203 797 2206
rect 818 2203 828 2206
rect 906 2203 940 2206
rect 1002 2203 1020 2206
rect 1300 2203 1309 2206
rect 1498 2203 1508 2206
rect 1556 2203 1565 2206
rect 1658 2203 1676 2206
rect 1698 2203 1732 2206
rect 1770 2203 1788 2206
rect 1866 2203 1869 2214
rect 1906 2213 1916 2216
rect 2028 2213 2061 2216
rect 2204 2213 2213 2216
rect 2226 2213 2244 2216
rect 2250 2213 2261 2216
rect 2292 2213 2316 2216
rect 2340 2213 2357 2216
rect 2258 2207 2261 2213
rect 2378 2207 2381 2216
rect 2444 2213 2460 2216
rect 2556 2213 2565 2216
rect 2066 2203 2076 2206
rect 2186 2203 2196 2206
rect 2308 2203 2317 2206
rect 2346 2203 2356 2206
rect 2386 2203 2395 2206
rect 2410 2203 2436 2206
rect 2578 2205 2581 2216
rect 2594 2213 2628 2216
rect 2586 2203 2604 2206
rect 2652 2203 2661 2206
rect 730 2193 772 2196
rect 818 2195 821 2203
rect 2410 2195 2413 2203
rect 2844 2176 2848 2472
rect -101 1876 -97 2172
rect 38 2167 2698 2173
rect 450 2136 453 2146
rect 2666 2136 2669 2156
rect 66 2133 76 2136
rect 212 2133 237 2136
rect 292 2133 325 2136
rect 450 2133 468 2136
rect 764 2133 773 2136
rect 812 2133 837 2136
rect 1164 2133 1172 2136
rect 1228 2133 1245 2136
rect 1260 2133 1277 2136
rect 1556 2133 1580 2136
rect 1596 2133 1613 2136
rect 1674 2133 1700 2136
rect 1740 2133 1757 2136
rect 84 2123 173 2126
rect 204 2123 213 2126
rect 244 2123 253 2126
rect 322 2123 325 2133
rect 450 2123 476 2126
rect 482 2123 492 2126
rect 714 2123 740 2126
rect 778 2123 796 2126
rect 884 2123 909 2126
rect 946 2123 964 2126
rect 1020 2123 1045 2126
rect 1180 2123 1189 2126
rect 1194 2123 1212 2126
rect 1234 2123 1252 2126
rect 1298 2123 1308 2126
rect 1234 2116 1237 2123
rect 1228 2113 1237 2116
rect 1474 2106 1477 2125
rect 1666 2123 1692 2126
rect 1724 2123 1732 2126
rect 1746 2123 1772 2126
rect 1802 2125 1805 2136
rect 1890 2125 1893 2136
rect 2098 2126 2101 2135
rect 2178 2133 2196 2136
rect 2244 2133 2261 2136
rect 2381 2133 2389 2136
rect 2410 2133 2420 2136
rect 2442 2126 2445 2135
rect 2610 2126 2613 2135
rect 2660 2133 2733 2136
rect 1956 2123 1989 2126
rect 2012 2123 2045 2126
rect 2068 2123 2101 2126
rect 2124 2123 2149 2126
rect 2204 2123 2228 2126
rect 2330 2123 2340 2126
rect 2346 2123 2364 2126
rect 2378 2123 2387 2126
rect 2436 2123 2445 2126
rect 2498 2123 2524 2126
rect 2546 2123 2580 2126
rect 2602 2123 2613 2126
rect 1778 2113 1788 2116
rect 1850 2113 1876 2116
rect 1890 2113 1900 2116
rect 2244 2113 2268 2116
rect 2292 2113 2300 2116
rect 682 2103 700 2106
rect 1466 2103 1477 2106
rect 2276 2103 2309 2106
rect 14 2067 2722 2073
rect 1524 2033 1541 2036
rect 642 2023 668 2026
rect 1484 2023 1493 2026
rect 1778 2016 1781 2025
rect 2252 2023 2261 2026
rect 2266 2016 2269 2025
rect 74 2013 84 2016
rect 210 2013 220 2016
rect 602 2013 612 2016
rect 698 2013 732 2016
rect 932 2013 957 2016
rect 1012 2013 1029 2016
rect 1042 2013 1052 2016
rect 1082 2013 1092 2016
rect 1132 2013 1181 2016
rect 1396 2013 1421 2016
rect 1452 2013 1461 2016
rect 1676 2013 1709 2016
rect 396 2003 429 2006
rect 434 2003 460 2006
rect 492 2003 501 2006
rect 698 2003 708 2006
rect 756 2003 773 2006
rect 1076 2003 1084 2006
rect 1098 2003 1108 2006
rect 1588 2003 1612 2006
rect 442 1993 445 2003
rect 1706 1996 1709 2013
rect 1730 2006 1733 2014
rect 1756 2013 1781 2016
rect 1730 2003 1748 2006
rect 1802 2003 1805 2014
rect 1836 2013 1885 2016
rect 2044 2013 2061 2016
rect 1866 2003 1900 2006
rect 1938 2003 1988 2006
rect 2068 2003 2109 2006
rect 2114 2003 2132 2006
rect 2146 2003 2149 2014
rect 2250 2013 2269 2016
rect 2276 2013 2293 2016
rect 2322 2013 2332 2016
rect 2364 2013 2380 2016
rect 2420 2013 2445 2016
rect 2452 2013 2476 2016
rect 2524 2013 2533 2016
rect 2546 2013 2557 2016
rect 2602 2013 2613 2016
rect 2636 2013 2645 2016
rect 2554 2005 2557 2013
rect 2610 2005 2613 2013
rect 2658 2006 2661 2016
rect 2658 2005 2669 2006
rect 2660 2003 2669 2005
rect 1698 1993 1716 1996
rect 2148 1993 2165 1996
rect 2316 1993 2325 1996
rect 38 1967 2698 1973
rect 514 1943 532 1946
rect 546 1936 549 1946
rect 1386 1936 1389 1945
rect 1818 1943 1844 1946
rect 2426 1943 2452 1946
rect 274 1933 292 1936
rect 308 1933 317 1936
rect 546 1933 556 1936
rect 570 1933 580 1936
rect 636 1933 661 1936
rect 780 1933 805 1936
rect 1362 1933 1372 1936
rect 1386 1933 1437 1936
rect 1482 1933 1492 1936
rect 252 1923 261 1926
rect 330 1923 348 1926
rect 554 1923 564 1926
rect 610 1923 620 1926
rect 676 1923 684 1926
rect 706 1923 740 1926
rect 834 1923 852 1926
rect 988 1923 997 1926
rect 1036 1923 1061 1926
rect 1124 1923 1149 1926
rect 1188 1923 1205 1926
rect 1284 1923 1309 1926
rect 1338 1923 1364 1926
rect 1434 1923 1437 1933
rect 1546 1926 1549 1935
rect 1610 1926 1613 1935
rect 1658 1933 1668 1936
rect 1690 1933 1708 1936
rect 1658 1926 1661 1933
rect 1458 1923 1500 1926
rect 1546 1923 1564 1926
rect 1602 1923 1613 1926
rect 1628 1923 1637 1926
rect 1652 1923 1661 1926
rect 1676 1923 1693 1926
rect 1738 1925 1741 1936
rect 1786 1933 1852 1936
rect 1882 1925 1885 1936
rect 1970 1923 1973 1935
rect 2074 1933 2092 1936
rect 2162 1933 2204 1936
rect 2284 1933 2293 1936
rect 2162 1925 2165 1933
rect 2370 1926 2373 1935
rect 2450 1933 2460 1936
rect 2212 1923 2229 1926
rect 2356 1923 2373 1926
rect 2394 1923 2412 1926
rect 2466 1925 2469 1946
rect 2530 1933 2540 1936
rect 2506 1923 2548 1926
rect 636 1913 645 1916
rect 834 1915 837 1923
rect 1756 1913 1781 1916
rect 2060 1913 2085 1916
rect 2250 1913 2260 1916
rect 2396 1913 2405 1916
rect 1882 1903 1892 1906
rect 2106 1903 2132 1906
rect 2844 1876 2848 2172
rect 14 1867 2722 1873
rect 412 1833 453 1836
rect 532 1833 549 1836
rect 722 1833 740 1836
rect 1396 1833 1413 1836
rect 1570 1833 1580 1836
rect 1882 1833 1901 1836
rect 2114 1833 2124 1836
rect 1882 1826 1885 1833
rect 148 1823 157 1826
rect 172 1823 189 1826
rect 298 1823 308 1826
rect 346 1823 356 1826
rect 394 1823 404 1826
rect 428 1823 445 1826
rect 500 1823 524 1826
rect 538 1823 548 1826
rect 748 1823 765 1826
rect 1370 1823 1388 1826
rect 1588 1823 1597 1826
rect 1868 1823 1885 1826
rect 1916 1823 1933 1826
rect 2482 1823 2524 1826
rect 146 1813 164 1816
rect 260 1813 277 1816
rect 90 1803 124 1806
rect 170 1803 188 1806
rect 202 1803 228 1806
rect 298 1803 301 1814
rect 324 1803 341 1806
rect 346 1796 349 1823
rect 460 1813 477 1816
rect 434 1803 452 1806
rect 474 1805 477 1813
rect 602 1813 620 1816
rect 500 1803 517 1806
rect 602 1805 605 1813
rect 642 1803 645 1814
rect 666 1806 669 1814
rect 700 1813 709 1816
rect 716 1813 732 1816
rect 828 1813 853 1816
rect 892 1813 917 1816
rect 956 1813 981 1816
rect 1058 1813 1076 1816
rect 1202 1813 1212 1816
rect 1308 1813 1341 1816
rect 1378 1806 1381 1823
rect 1666 1813 1692 1816
rect 1748 1813 1772 1816
rect 1794 1813 1813 1816
rect 1972 1813 2005 1816
rect 2058 1813 2084 1816
rect 666 1803 677 1806
rect 754 1803 772 1806
rect 786 1803 820 1806
rect 834 1803 860 1806
rect 1028 1803 1045 1806
rect 1084 1803 1101 1806
rect 1146 1803 1204 1806
rect 1316 1803 1381 1806
rect 1434 1803 1444 1806
rect 1514 1803 1540 1806
rect 1668 1803 1677 1806
rect 1682 1803 1724 1806
rect 1740 1803 1749 1806
rect 1786 1803 1796 1806
rect 1810 1805 1813 1813
rect 2002 1806 2005 1813
rect 2002 1803 2028 1806
rect 2044 1803 2069 1806
rect 2114 1803 2117 1814
rect 2156 1813 2165 1816
rect 2186 1813 2204 1816
rect 2258 1813 2268 1816
rect 2138 1803 2148 1806
rect 2154 1803 2164 1806
rect 2298 1803 2316 1806
rect 2362 1803 2365 1814
rect 2418 1813 2445 1816
rect 2476 1813 2485 1816
rect 2420 1803 2429 1806
rect 2444 1803 2460 1806
rect 2562 1803 2565 1814
rect 2626 1813 2644 1816
rect 2602 1803 2612 1806
rect 2618 1803 2636 1806
rect 332 1793 349 1796
rect 1514 1793 1532 1796
rect 2292 1793 2308 1796
rect 38 1767 2698 1773
rect 74 1743 92 1746
rect 332 1743 364 1746
rect 514 1743 532 1746
rect 586 1743 612 1746
rect 106 1733 124 1736
rect 108 1723 125 1726
rect 132 1723 157 1726
rect 162 1725 165 1736
rect 244 1733 277 1736
rect 346 1733 372 1736
rect 378 1733 396 1736
rect 450 1726 453 1735
rect 476 1733 485 1736
rect 500 1733 533 1736
rect 540 1733 557 1736
rect 610 1733 620 1736
rect 178 1723 196 1726
rect 380 1723 389 1726
rect 428 1723 453 1726
rect 474 1723 492 1726
rect 554 1725 557 1733
rect 580 1723 613 1726
rect 626 1725 629 1736
rect 642 1725 645 1736
rect 730 1726 733 1735
rect 802 1726 805 1735
rect 908 1733 925 1736
rect 1002 1733 1036 1736
rect 722 1723 733 1726
rect 794 1723 805 1726
rect 836 1723 861 1726
rect 892 1723 941 1726
rect 978 1723 1028 1726
rect 1058 1725 1061 1736
rect 1074 1733 1092 1736
rect 1114 1733 1140 1736
rect 1066 1723 1084 1726
rect 1122 1723 1132 1726
rect 1180 1723 1197 1726
rect 1298 1725 1301 1736
rect 1308 1733 1317 1736
rect 1332 1733 1348 1736
rect 1370 1733 1380 1736
rect 1324 1723 1333 1726
rect 1370 1725 1373 1733
rect 1434 1726 1437 1735
rect 1458 1726 1461 1735
rect 1532 1733 1549 1736
rect 1586 1733 1596 1736
rect 1706 1726 1709 1735
rect 1762 1726 1765 1735
rect 1818 1726 1821 1735
rect 1922 1726 1925 1735
rect 1930 1733 1940 1736
rect 1988 1733 1997 1736
rect 1404 1723 1437 1726
rect 1444 1723 1461 1726
rect 1610 1723 1620 1726
rect 1676 1723 1709 1726
rect 1738 1723 1765 1726
rect 1794 1723 1821 1726
rect 1906 1723 1925 1726
rect 2002 1726 2005 1735
rect 2074 1733 2116 1736
rect 2002 1723 2021 1726
rect 2146 1725 2149 1736
rect 2386 1733 2428 1736
rect 2322 1723 2348 1726
rect 2354 1723 2364 1726
rect 2474 1725 2477 1736
rect 2490 1725 2493 1746
rect 2508 1743 2525 1746
rect 2546 1733 2556 1736
rect 2562 1726 2565 1745
rect 2506 1723 2532 1726
rect 2538 1723 2548 1726
rect 2562 1723 2573 1726
rect 2634 1725 2637 1736
rect 722 1716 725 1723
rect 794 1716 797 1723
rect 674 1713 684 1716
rect 708 1713 725 1716
rect 746 1713 756 1716
rect 780 1713 797 1716
rect 2186 1713 2196 1716
rect 2570 1715 2573 1723
rect 2602 1713 2620 1716
rect 2634 1713 2644 1716
rect 634 1703 652 1706
rect 666 1703 700 1706
rect 1482 1703 1492 1706
rect 2138 1703 2156 1706
rect 14 1667 2722 1673
rect 130 1633 188 1636
rect 330 1633 340 1636
rect 1420 1633 1453 1636
rect 1522 1633 1548 1636
rect 2388 1633 2397 1636
rect 138 1623 172 1626
rect 260 1623 269 1626
rect 348 1623 365 1626
rect 1402 1623 1412 1626
rect 1426 1623 1436 1626
rect 1514 1623 1532 1626
rect 2434 1623 2444 1626
rect 124 1613 165 1616
rect 316 1613 332 1616
rect 412 1613 421 1616
rect 444 1613 452 1616
rect 524 1613 573 1616
rect 676 1613 725 1616
rect 354 1603 372 1606
rect 474 1603 492 1606
rect 554 1603 572 1606
rect 636 1603 645 1606
rect 842 1603 845 1614
rect 876 1613 885 1616
rect 874 1603 884 1606
rect 994 1603 997 1614
rect 1034 1613 1084 1616
rect 1106 1613 1148 1616
rect 1178 1606 1181 1614
rect 1186 1613 1228 1616
rect 1298 1613 1325 1616
rect 1332 1613 1373 1616
rect 1020 1603 1029 1606
rect 1042 1603 1060 1606
rect 1138 1603 1156 1606
rect 1178 1603 1204 1606
rect 1292 1603 1301 1606
rect 1322 1605 1325 1613
rect 1402 1606 1405 1623
rect 1442 1613 1460 1616
rect 1562 1613 1580 1616
rect 1618 1613 1644 1616
rect 1674 1613 1700 1616
rect 1756 1613 1765 1616
rect 1818 1613 1845 1616
rect 2018 1613 2037 1616
rect 2266 1613 2285 1616
rect 2308 1613 2333 1616
rect 1388 1603 1405 1606
rect 1450 1603 1468 1606
rect 1482 1603 1509 1606
rect 1724 1603 1732 1606
rect 1842 1605 1845 1613
rect 1892 1603 1917 1606
rect 2018 1603 2036 1606
rect 2084 1603 2109 1606
rect 2164 1603 2173 1606
rect 2178 1603 2204 1606
rect 2252 1603 2277 1606
rect 2332 1603 2341 1606
rect 2484 1603 2501 1606
rect 2530 1603 2533 1614
rect 2546 1603 2556 1606
rect 2660 1603 2669 1606
rect 1482 1597 1485 1603
rect 124 1593 149 1596
rect 1508 1593 1517 1596
rect 2844 1576 2848 1872
rect 38 1567 2698 1573
rect 1298 1536 1301 1545
rect 706 1526 709 1535
rect 714 1533 724 1536
rect 386 1523 396 1526
rect 426 1523 452 1526
rect 524 1523 549 1526
rect 580 1523 605 1526
rect 636 1523 661 1526
rect 690 1523 716 1526
rect 746 1525 749 1536
rect 842 1533 852 1536
rect 978 1533 988 1536
rect 1010 1533 1044 1536
rect 1260 1533 1268 1536
rect 1292 1533 1301 1536
rect 780 1523 812 1526
rect 844 1523 853 1526
rect 1012 1523 1029 1526
rect 1202 1523 1236 1526
rect 1284 1523 1301 1526
rect 1314 1525 1317 1536
rect 1338 1533 1348 1536
rect 1370 1533 1388 1536
rect 1402 1533 1412 1536
rect 1434 1533 1460 1536
rect 1476 1533 1485 1536
rect 1556 1533 1565 1536
rect 1596 1526 1613 1527
rect 1658 1526 1661 1535
rect 1778 1526 1781 1535
rect 1898 1533 1916 1536
rect 1980 1533 1997 1536
rect 2052 1533 2085 1536
rect 2140 1533 2149 1536
rect 2372 1533 2389 1536
rect 2490 1533 2508 1536
rect 2546 1533 2572 1536
rect 2596 1533 2605 1536
rect 2660 1533 2733 1536
rect 1372 1523 1381 1526
rect 1436 1523 1452 1526
rect 1522 1523 1532 1526
rect 1538 1523 1548 1526
rect 1596 1524 1628 1526
rect 1610 1523 1628 1524
rect 1658 1523 1692 1526
rect 1748 1523 1781 1526
rect 2002 1523 2020 1526
rect 2226 1523 2236 1526
rect 2276 1523 2325 1526
rect 2354 1523 2364 1526
rect 292 1513 300 1516
rect 1026 1513 1029 1523
rect 1538 1515 1541 1523
rect 1570 1513 1580 1516
rect 1594 1513 1604 1516
rect 2378 1513 2396 1516
rect 2442 1513 2452 1516
rect 2490 1506 2493 1533
rect 2514 1523 2524 1526
rect 2548 1523 2565 1526
rect 2594 1523 2636 1526
rect 276 1503 316 1506
rect 330 1503 348 1506
rect 1588 1503 1605 1506
rect 2436 1503 2453 1506
rect 2474 1503 2493 1506
rect 14 1472 2722 1473
rect 6 1468 2722 1472
rect 6 1452 10 1468
rect 14 1467 2722 1468
rect -117 1448 10 1452
rect -102 1276 -98 1448
rect 1396 1433 1421 1436
rect 124 1423 133 1426
rect 1316 1423 1324 1426
rect 1362 1423 1388 1426
rect 2482 1423 2492 1426
rect 2578 1416 2581 1425
rect 154 1413 164 1416
rect 180 1403 205 1406
rect 266 1403 269 1414
rect 284 1413 293 1416
rect 324 1413 341 1416
rect 306 1403 316 1406
rect 394 1403 397 1414
rect 524 1413 565 1416
rect 596 1413 629 1416
rect 668 1413 693 1416
rect 724 1413 741 1416
rect 788 1413 797 1416
rect 850 1413 884 1416
rect 922 1413 932 1416
rect 1050 1413 1060 1416
rect 1116 1413 1141 1416
rect 1146 1413 1172 1416
rect 1194 1413 1204 1416
rect 1236 1413 1261 1416
rect 1266 1413 1276 1416
rect 1466 1413 1476 1416
rect 1498 1413 1508 1416
rect 1540 1413 1548 1416
rect 1562 1413 1580 1416
rect 1604 1413 1613 1416
rect 1628 1413 1653 1416
rect 1916 1413 1949 1416
rect 2002 1413 2020 1416
rect 2252 1413 2261 1416
rect 2468 1413 2477 1416
rect 2508 1413 2533 1416
rect 2546 1413 2556 1416
rect 2562 1413 2581 1416
rect 450 1403 484 1406
rect 548 1403 557 1406
rect 620 1403 637 1406
rect 692 1403 701 1406
rect 738 1405 741 1413
rect 754 1403 764 1406
rect 786 1403 836 1406
rect 850 1403 892 1406
rect 914 1403 924 1406
rect 1196 1403 1205 1406
rect 1234 1403 1268 1406
rect 1418 1403 1428 1406
rect 1490 1403 1516 1406
rect 1556 1403 1573 1406
rect 1602 1403 1620 1406
rect 1858 1403 1892 1406
rect 1908 1403 2028 1406
rect 2050 1403 2060 1406
rect 2386 1403 2396 1406
rect 2466 1403 2492 1406
rect 2522 1403 2548 1406
rect 218 1393 252 1396
rect 2434 1393 2444 1396
rect 38 1367 2698 1373
rect 106 1343 116 1346
rect 1458 1343 1484 1346
rect 2380 1343 2389 1346
rect 2458 1343 2468 1346
rect 98 1323 116 1326
rect 154 1323 164 1326
rect 306 1325 309 1336
rect 322 1325 325 1336
rect 346 1333 372 1336
rect 706 1333 748 1336
rect 1044 1333 1069 1336
rect 1074 1333 1108 1336
rect 1130 1333 1180 1336
rect 1428 1333 1437 1336
rect 1442 1326 1445 1335
rect 1458 1333 1492 1336
rect 354 1323 380 1326
rect 426 1323 436 1326
rect 690 1323 740 1326
rect 842 1323 852 1326
rect 1052 1323 1061 1326
rect 1082 1323 1100 1326
rect 1132 1323 1149 1326
rect 1154 1323 1172 1326
rect 1204 1323 1213 1326
rect 1260 1323 1269 1326
rect 1322 1323 1348 1326
rect 1402 1323 1413 1326
rect 1420 1323 1445 1326
rect 1452 1323 1485 1326
rect 1498 1325 1501 1336
rect 1516 1333 1548 1336
rect 1780 1333 1797 1336
rect 1826 1333 1876 1336
rect 1898 1333 1908 1336
rect 2346 1326 2349 1335
rect 2372 1333 2381 1336
rect 2436 1333 2452 1336
rect 2514 1333 2524 1336
rect 1514 1323 1540 1326
rect 1572 1323 1580 1326
rect 1618 1323 1628 1326
rect 1634 1323 1644 1326
rect 1778 1323 1796 1326
rect 1828 1323 1861 1326
rect 2066 1323 2092 1326
rect 2298 1323 2316 1326
rect 2346 1323 2356 1326
rect 2412 1324 2428 1327
rect 2546 1326 2549 1335
rect 2570 1333 2580 1336
rect 2492 1323 2501 1326
rect 2508 1323 2525 1326
rect 2546 1323 2564 1326
rect 2578 1323 2596 1326
rect 340 1313 365 1316
rect 492 1313 501 1316
rect 522 1313 532 1316
rect 570 1313 588 1316
rect 1402 1315 1405 1323
rect 1634 1315 1637 1323
rect 2386 1313 2396 1316
rect 314 1303 332 1306
rect 474 1303 484 1306
rect 2404 1303 2413 1306
rect 2844 1276 2848 1572
rect -102 976 -98 1272
rect 14 1267 2722 1273
rect 130 1233 148 1236
rect 1458 1233 1484 1236
rect 2530 1233 2548 1236
rect 132 1223 141 1226
rect 1492 1223 1501 1226
rect 114 1213 124 1216
rect 162 1213 172 1216
rect 316 1213 325 1216
rect 330 1213 357 1216
rect 388 1213 413 1216
rect 428 1213 437 1216
rect 484 1213 517 1216
rect 556 1213 564 1216
rect 106 1203 116 1206
rect 354 1196 357 1213
rect 490 1203 532 1206
rect 548 1203 565 1206
rect 594 1203 597 1214
rect 650 1213 684 1216
rect 794 1213 820 1216
rect 906 1213 917 1216
rect 906 1205 909 1213
rect 914 1205 917 1213
rect 962 1205 965 1216
rect 1098 1213 1117 1216
rect 1114 1205 1117 1213
rect 1122 1205 1125 1216
rect 1234 1205 1237 1216
rect 1346 1213 1372 1216
rect 1434 1213 1453 1216
rect 1458 1213 1476 1216
rect 1546 1213 1596 1216
rect 1746 1213 1772 1216
rect 1804 1213 1813 1216
rect 1450 1206 1453 1213
rect 1450 1205 1461 1206
rect 1452 1203 1461 1205
rect 1546 1203 1549 1213
rect 1612 1203 1621 1206
rect 1740 1203 1773 1206
rect 1858 1205 1861 1216
rect 1874 1213 1900 1216
rect 1930 1213 1956 1216
rect 1994 1213 2012 1216
rect 2044 1213 2069 1216
rect 2172 1213 2285 1216
rect 2308 1213 2341 1216
rect 2346 1213 2364 1216
rect 2412 1213 2429 1216
rect 1988 1203 2013 1206
rect 2036 1203 2061 1206
rect 2066 1205 2069 1213
rect 2116 1203 2141 1206
rect 2274 1203 2284 1206
rect 2338 1203 2341 1213
rect 2378 1203 2396 1206
rect 2420 1203 2429 1206
rect 2434 1203 2437 1214
rect 2468 1213 2476 1216
rect 2460 1203 2469 1206
rect 2522 1203 2525 1214
rect 2562 1213 2580 1216
rect 2602 1206 2605 1214
rect 2618 1213 2636 1216
rect 2602 1203 2644 1206
rect 354 1193 364 1196
rect 1530 1193 1565 1196
rect 1620 1193 1629 1196
rect 2498 1193 2508 1196
rect 38 1167 2698 1173
rect 1034 1153 1061 1156
rect 538 1143 548 1146
rect 1034 1143 1053 1146
rect 170 1126 173 1135
rect 452 1133 477 1136
rect 498 1133 508 1136
rect 530 1133 556 1136
rect 604 1133 613 1136
rect 660 1133 684 1136
rect 868 1133 885 1136
rect 890 1126 893 1135
rect 940 1133 965 1136
rect 970 1133 980 1136
rect 1028 1133 1053 1136
rect 1108 1133 1125 1136
rect 1162 1133 1180 1136
rect 1194 1126 1197 1135
rect 1210 1133 1388 1136
rect 1434 1126 1437 1135
rect 1780 1133 1813 1136
rect 1842 1133 1852 1136
rect 108 1123 133 1126
rect 164 1123 173 1126
rect 466 1123 484 1126
rect 532 1123 541 1126
rect 570 1123 596 1126
rect 666 1123 700 1126
rect 762 1123 788 1126
rect 874 1123 893 1126
rect 938 1123 1004 1126
rect 1114 1123 1197 1126
rect 1370 1123 1412 1126
rect 1434 1123 1445 1126
rect 1588 1123 1621 1126
rect 1708 1123 1733 1126
rect 1794 1123 1812 1126
rect 1844 1123 1853 1126
rect 1986 1123 1996 1126
rect 2018 1123 2044 1126
rect 2138 1125 2141 1136
rect 2170 1133 2180 1136
rect 2290 1126 2293 1135
rect 2284 1123 2293 1126
rect 2402 1125 2405 1136
rect 2452 1133 2485 1136
rect 2522 1126 2525 1135
rect 2634 1133 2644 1136
rect 2426 1123 2444 1126
rect 2522 1123 2533 1126
rect 1442 1116 1445 1123
rect 2530 1116 2533 1123
rect 610 1113 620 1116
rect 1442 1113 1476 1116
rect 1506 1113 1532 1116
rect 2386 1113 2396 1116
rect 2420 1113 2437 1116
rect 2530 1113 2540 1116
rect 1484 1103 1525 1106
rect 2364 1103 2373 1106
rect 2386 1093 2389 1113
rect 2612 1103 2621 1106
rect 14 1067 2722 1073
rect 2340 1033 2357 1036
rect 2468 1033 2509 1036
rect 300 1023 309 1026
rect 322 1016 325 1025
rect 698 1023 708 1026
rect 2322 1023 2332 1026
rect 2474 1023 2484 1026
rect 2322 1016 2325 1023
rect 58 1013 69 1016
rect 108 1013 133 1016
rect 146 1013 156 1016
rect 188 1013 197 1016
rect 58 996 61 1013
rect 66 1003 76 1006
rect 194 1005 197 1013
rect 226 1003 229 1014
rect 322 1013 332 1016
rect 354 1013 364 1016
rect 370 1013 381 1016
rect 426 1013 444 1016
rect 474 1013 493 1016
rect 522 1013 540 1016
rect 602 1013 612 1016
rect 340 1003 349 1006
rect 370 1005 373 1013
rect 474 1005 477 1013
rect 524 1003 533 1006
rect 562 1003 580 1006
rect 602 1005 605 1013
rect 658 1006 661 1014
rect 698 1013 716 1016
rect 722 1013 756 1016
rect 786 1013 804 1016
rect 874 1013 924 1016
rect 946 1013 956 1016
rect 698 1006 701 1013
rect 644 1003 661 1006
rect 684 1003 709 1006
rect 722 1005 725 1013
rect 1098 1006 1101 1016
rect 1148 1013 1165 1016
rect 1204 1013 1244 1016
rect 1274 1006 1277 1014
rect 1420 1013 1453 1016
rect 1476 1013 1485 1016
rect 1618 1013 1637 1016
rect 1764 1013 1789 1016
rect 1826 1013 1844 1016
rect 1850 1013 1876 1016
rect 1908 1013 1949 1016
rect 2010 1013 2060 1016
rect 2090 1013 2100 1016
rect 2244 1013 2253 1016
rect 2266 1013 2276 1016
rect 2298 1013 2308 1016
rect 2314 1013 2325 1016
rect 1050 1003 1060 1006
rect 1084 1003 1093 1006
rect 1098 1003 1140 1006
rect 1146 1003 1196 1006
rect 1274 1003 1285 1006
rect 1306 1003 1324 1006
rect 1330 1003 1340 1006
rect 1450 1005 1453 1013
rect 1618 1005 1621 1013
rect 2010 1006 2013 1013
rect 1852 1003 1877 1006
rect 1930 1003 1948 1006
rect 1996 1003 2013 1006
rect 2018 1003 2044 1006
rect 2092 1003 2101 1006
rect 2130 1003 2140 1006
rect 2250 1005 2253 1013
rect 2314 1005 2317 1013
rect 2394 1006 2397 1014
rect 2372 1003 2381 1006
rect 2394 1003 2428 1006
rect 2474 1003 2477 1014
rect 2618 1013 2636 1016
rect 2498 1003 2524 1006
rect 2538 1003 2564 1006
rect 2604 1003 2629 1006
rect 2644 1003 2709 1006
rect 1090 996 1093 1003
rect 58 993 69 996
rect 626 993 636 996
rect 1090 993 1132 996
rect 1282 995 1285 1003
rect 2378 995 2381 1003
rect 2532 993 2557 996
rect 66 983 69 993
rect -102 676 -98 972
rect 38 967 2698 973
rect 580 943 589 946
rect 658 943 668 946
rect 1268 943 1277 946
rect 2258 943 2277 946
rect 2274 936 2277 943
rect 2706 936 2709 1003
rect 108 923 125 926
rect 290 923 293 934
rect 314 925 317 936
rect 338 925 341 936
rect 402 925 405 936
rect 492 933 517 936
rect 556 933 565 936
rect 690 933 701 936
rect 458 923 468 926
rect 506 923 532 926
rect 626 923 668 926
rect 690 925 693 933
rect 698 923 716 926
rect 722 923 748 926
rect 810 925 813 936
rect 948 933 957 936
rect 1066 926 1069 934
rect 842 923 868 926
rect 914 923 924 926
rect 946 923 965 926
rect 1058 923 1069 926
rect 1076 923 1092 926
rect 1122 925 1125 936
rect 1154 925 1157 936
rect 1178 933 1212 936
rect 1234 925 1237 936
rect 1260 933 1277 936
rect 1274 926 1277 933
rect 1274 923 1300 926
rect 1306 923 1324 926
rect 1354 925 1357 936
rect 1420 933 1428 936
rect 1474 926 1477 934
rect 1386 923 1396 926
rect 1474 923 1485 926
rect 1586 923 1589 934
rect 1594 923 1597 934
rect 1818 933 1844 936
rect 1892 933 1909 936
rect 1930 933 1940 936
rect 1988 933 1997 936
rect 2066 933 2140 936
rect 2170 933 2188 936
rect 2252 933 2269 936
rect 2274 933 2284 936
rect 2298 933 2316 936
rect 1642 923 1676 926
rect 2036 923 2125 926
rect 2164 923 2189 926
rect 2282 923 2292 926
rect 2378 925 2381 936
rect 2396 933 2413 936
rect 2404 923 2452 926
rect 2482 923 2485 934
rect 2538 925 2541 936
rect 2570 925 2573 936
rect 2610 926 2613 934
rect 2660 933 2709 936
rect 2602 923 2613 926
rect 1058 916 1061 923
rect 292 913 300 916
rect 356 913 365 916
rect 420 913 429 916
rect 586 913 596 916
rect 778 913 796 916
rect 810 913 820 916
rect 1036 913 1061 916
rect 1130 913 1148 916
rect 1306 915 1309 923
rect 1354 913 1364 916
rect 308 903 341 906
rect 394 903 412 906
rect 426 893 429 913
rect 586 903 612 906
rect 988 903 997 906
rect 1020 903 1061 906
rect 1146 903 1164 906
rect 2498 903 2524 906
rect 14 867 2722 873
rect 2845 848 2865 852
rect 1500 833 1509 836
rect 2226 833 2252 836
rect 194 816 197 825
rect 906 823 916 826
rect 1482 823 1492 826
rect 2236 823 2245 826
rect 2260 823 2277 826
rect 2314 823 2332 826
rect 2484 823 2501 826
rect 2498 816 2501 823
rect 180 813 197 816
rect 260 813 285 816
rect 322 813 332 816
rect 186 803 196 806
rect 386 805 389 816
rect 492 813 509 816
rect 516 813 565 816
rect 612 813 637 816
rect 660 813 669 816
rect 506 805 509 813
rect 570 803 588 806
rect 604 803 613 806
rect 642 803 652 806
rect 682 803 685 814
rect 754 813 788 816
rect 876 813 901 816
rect 986 813 1004 816
rect 1074 813 1092 816
rect 1074 806 1077 813
rect 812 803 820 806
rect 844 803 861 806
rect 1060 803 1077 806
rect 1106 805 1109 816
rect 1116 813 1125 816
rect 1170 813 1204 816
rect 1226 813 1237 816
rect 1170 805 1173 813
rect 1226 805 1229 813
rect 1234 805 1237 813
rect 1282 813 1316 816
rect 1372 813 1405 816
rect 1418 813 1452 816
rect 1610 813 1620 816
rect 1282 805 1285 813
rect 1476 803 1485 806
rect 1522 803 1532 806
rect 1642 803 1668 806
rect 1722 805 1725 816
rect 1748 813 1757 816
rect 1874 813 1916 816
rect 1954 813 1980 816
rect 2012 813 2021 816
rect 1826 803 1844 806
rect 1866 803 1924 806
rect 1946 803 1988 806
rect 2010 803 2020 806
rect 2034 803 2044 806
rect 2090 805 2093 816
rect 2106 805 2109 816
rect 2162 813 2205 816
rect 2162 806 2165 813
rect 2148 803 2165 806
rect 1644 793 1661 796
rect 2202 795 2205 813
rect 2212 803 2229 806
rect 2242 803 2245 814
rect 2266 813 2284 816
rect 2386 813 2404 816
rect 2458 813 2476 816
rect 2498 813 2565 816
rect 2572 813 2589 816
rect 2602 813 2636 816
rect 2314 803 2332 806
rect 2386 805 2389 813
rect 2426 803 2436 806
rect 2458 805 2461 813
rect 2506 803 2516 806
rect 2538 803 2564 806
rect 2658 805 2661 816
rect 2314 796 2317 803
rect 2308 793 2317 796
rect 38 767 2698 773
rect 2284 743 2293 746
rect 186 733 196 736
rect 236 733 261 736
rect 284 733 317 736
rect 322 726 325 735
rect 354 733 388 736
rect 442 733 468 736
rect 570 726 573 735
rect 180 723 197 726
rect 212 723 269 726
rect 276 723 325 726
rect 508 723 541 726
rect 570 723 581 726
rect 602 725 605 736
rect 660 733 677 736
rect 740 733 749 736
rect 844 733 853 736
rect 924 733 956 736
rect 642 723 652 726
rect 836 723 869 726
rect 922 723 948 726
rect 980 723 989 726
rect 1042 725 1045 736
rect 1108 733 1125 736
rect 1364 733 1372 736
rect 1476 733 1493 736
rect 1498 726 1501 735
rect 1554 733 1572 736
rect 1058 723 1100 726
rect 1138 723 1172 726
rect 1402 723 1452 726
rect 1474 723 1501 726
rect 1538 723 1548 726
rect 1596 723 1605 726
rect 1690 723 1716 726
rect 1786 723 1796 726
rect 1842 723 1852 726
rect 1946 723 1956 726
rect 2162 723 2173 726
rect 2186 725 2189 736
rect 2266 733 2276 736
rect 2282 733 2308 736
rect 2394 733 2420 736
rect 2652 733 2669 736
rect 2282 723 2316 726
rect 2332 723 2341 726
rect 2428 723 2437 726
rect 2530 723 2556 726
rect 2596 723 2605 726
rect 2618 723 2628 726
rect 194 715 197 723
rect 578 716 581 723
rect 348 713 381 716
rect 578 713 588 716
rect 612 713 621 716
rect 866 706 869 723
rect 2170 716 2173 723
rect 900 713 909 716
rect 986 713 1028 716
rect 1042 713 1052 716
rect 1610 713 1660 716
rect 2170 713 2180 716
rect 2218 713 2236 716
rect 2340 713 2349 716
rect 2500 713 2509 716
rect 866 703 892 706
rect 2210 703 2252 706
rect 2845 677 2849 848
rect -102 376 -98 672
rect 14 667 2722 673
rect 2436 633 2469 636
rect 2154 623 2196 626
rect 2418 623 2428 626
rect 204 613 229 616
rect 412 613 445 616
rect 628 613 645 616
rect 706 613 732 616
rect 850 613 860 616
rect 964 613 972 616
rect 978 613 988 616
rect 1012 613 1021 616
rect 1116 613 1140 616
rect 1210 613 1220 616
rect 1244 613 1253 616
rect 1266 613 1324 616
rect 1362 613 1396 616
rect 1436 613 1453 616
rect 1468 613 1477 616
rect 1546 613 1556 616
rect 1580 613 1589 616
rect 1604 613 1612 616
rect 442 605 445 613
rect 642 605 645 613
rect 906 603 940 606
rect 980 603 989 606
rect 1010 603 1028 606
rect 1092 603 1101 606
rect 1164 603 1196 606
rect 1250 605 1253 613
rect 1298 603 1308 606
rect 1442 603 1452 606
rect 1562 603 1572 606
rect 1610 603 1620 606
rect 1642 603 1645 614
rect 1658 613 1668 616
rect 1690 603 1708 606
rect 1714 603 1717 614
rect 1722 613 1748 616
rect 1874 613 1893 616
rect 1930 613 1964 616
rect 2042 613 2076 616
rect 2140 613 2173 616
rect 2212 613 2237 616
rect 1874 605 1877 613
rect 1988 603 1996 606
rect 2042 605 2045 613
rect 2242 606 2245 614
rect 2306 613 2316 616
rect 2354 613 2380 616
rect 2092 603 2124 606
rect 2148 603 2165 606
rect 2178 603 2196 606
rect 2220 603 2245 606
rect 2266 603 2308 606
rect 2322 603 2364 606
rect 2442 603 2445 614
rect 2458 613 2484 616
rect 2516 613 2525 616
rect 2530 603 2533 614
rect 2556 603 2565 606
rect 2570 603 2573 614
rect 2620 613 2637 616
rect 2594 603 2612 606
rect 2618 603 2636 606
rect 1204 593 1213 596
rect 2100 593 2109 596
rect 2266 595 2269 603
rect 38 567 2698 573
rect 1410 536 1413 545
rect 202 533 212 536
rect 258 526 261 535
rect 386 526 389 535
rect 690 533 708 536
rect 196 523 213 526
rect 228 523 261 526
rect 324 523 341 526
rect 380 523 389 526
rect 572 523 597 526
rect 676 523 693 526
rect 754 525 757 536
rect 794 525 797 536
rect 826 533 844 536
rect 874 526 877 535
rect 986 526 989 535
rect 1330 533 1348 536
rect 868 523 893 526
rect 986 523 1005 526
rect 1196 523 1213 526
rect 1266 523 1276 526
rect 1282 523 1292 526
rect 1298 523 1308 526
rect 1332 523 1341 526
rect 1354 525 1357 536
rect 1404 533 1413 536
rect 1434 533 1444 536
rect 1572 533 1581 536
rect 1610 526 1613 545
rect 2274 543 2356 546
rect 2418 543 2444 546
rect 2572 543 2581 546
rect 2578 536 2581 543
rect 1676 533 1693 536
rect 1748 533 1789 536
rect 1956 533 2013 536
rect 2068 533 2101 536
rect 1460 523 1469 526
rect 1530 523 1548 526
rect 1586 523 1613 526
rect 1634 523 1652 526
rect 1714 523 1724 526
rect 1810 523 1820 526
rect 1850 523 1876 526
rect 1898 523 1932 526
rect 1954 523 2044 526
rect 2314 523 2356 526
rect 2378 525 2381 536
rect 2412 523 2421 526
rect 2442 525 2445 536
rect 2506 533 2516 536
rect 2570 533 2596 536
rect 2522 523 2556 526
rect 210 515 213 523
rect 660 513 669 516
rect 684 513 693 516
rect 1124 513 1133 516
rect 1210 513 1220 516
rect 1282 515 1285 523
rect 1514 513 1524 516
rect 2148 513 2181 516
rect 2186 513 2236 516
rect 2260 513 2269 516
rect 2314 513 2317 523
rect 690 503 693 513
rect 1108 503 1125 506
rect 2244 503 2301 506
rect 2484 503 2493 506
rect 14 467 2722 473
rect 1348 433 1365 436
rect 1602 433 1612 436
rect 1852 433 1861 436
rect 2404 433 2413 436
rect 194 416 197 425
rect 1082 423 1108 426
rect 1306 423 1340 426
rect 2386 423 2396 426
rect 2410 423 2420 426
rect 2588 423 2596 426
rect 66 413 76 416
rect 180 413 197 416
rect 212 413 221 416
rect 378 413 388 416
rect 186 403 196 406
rect 562 403 565 414
rect 594 403 597 414
rect 652 413 677 416
rect 732 413 741 416
rect 940 413 965 416
rect 970 413 980 416
rect 1018 413 1052 416
rect 1252 413 1268 416
rect 1300 413 1317 416
rect 1500 413 1509 416
rect 1540 413 1565 416
rect 1642 413 1756 416
rect 932 403 988 406
rect 1076 403 1101 406
rect 1156 403 1165 406
rect 1170 403 1188 406
rect 1244 403 1253 406
rect 1266 403 1276 406
rect 1386 403 1420 406
rect 1482 403 1492 406
rect 1498 403 1508 406
rect 1674 403 1732 406
rect 1778 405 1781 416
rect 1786 413 1812 416
rect 1860 413 1876 416
rect 1882 413 1924 416
rect 2010 406 2013 414
rect 2106 413 2156 416
rect 2330 413 2356 416
rect 2476 413 2500 416
rect 2524 413 2541 416
rect 2548 413 2557 416
rect 2612 413 2644 416
rect 1884 403 1893 406
rect 2010 403 2028 406
rect 2506 403 2516 406
rect 2538 405 2541 413
rect 2626 403 2636 406
rect 1164 393 1181 396
rect 2380 393 2389 396
rect 2845 376 2849 673
rect -102 76 -98 372
rect 38 367 2698 373
rect 1426 343 1476 346
rect 1602 336 1605 346
rect 1812 343 1821 346
rect 2578 336 2581 345
rect 186 333 196 336
rect 226 333 260 336
rect 274 326 277 335
rect 306 333 316 336
rect 356 333 373 336
rect 388 333 413 336
rect 426 333 436 336
rect 490 333 540 336
rect 666 326 669 335
rect 682 333 692 336
rect 716 333 741 336
rect 882 326 885 335
rect 948 333 981 336
rect 1010 333 1036 336
rect 1058 333 1068 336
rect 1122 333 1140 336
rect 1188 333 1205 336
rect 1316 333 1349 336
rect 1492 333 1548 336
rect 1570 326 1573 335
rect 1602 333 1620 336
rect 1682 333 1692 336
rect 1804 333 1813 336
rect 1890 326 1893 335
rect 66 323 76 326
rect 180 323 197 326
rect 212 323 261 326
rect 268 323 277 326
rect 314 323 324 326
rect 330 323 348 326
rect 380 323 421 326
rect 434 323 444 326
rect 522 323 532 326
rect 604 323 629 326
rect 660 323 669 326
rect 676 323 693 326
rect 708 323 717 326
rect 820 323 845 326
rect 876 323 885 326
rect 898 323 924 326
rect 1060 323 1085 326
rect 1130 323 1164 326
rect 1426 323 1476 326
rect 1500 323 1549 326
rect 1556 323 1573 326
rect 1602 323 1637 326
rect 1644 323 1653 326
rect 1770 323 1788 326
rect 1882 323 1893 326
rect 1914 326 1917 335
rect 1946 333 1957 336
rect 2026 333 2036 336
rect 1914 323 1924 326
rect 1946 325 1949 333
rect 2068 323 2085 326
rect 2092 323 2100 326
rect 2130 325 2133 336
rect 2204 333 2220 336
rect 2324 333 2333 336
rect 2138 323 2188 326
rect 2236 323 2253 326
rect 2338 323 2356 326
rect 2394 325 2397 336
rect 2410 325 2413 336
rect 2450 333 2468 336
rect 2482 333 2492 336
rect 2546 326 2549 335
rect 2572 333 2581 336
rect 2602 333 2612 336
rect 2476 323 2493 326
rect 2532 323 2549 326
rect 2604 323 2628 326
rect 194 315 197 323
rect 300 313 309 316
rect 460 313 501 316
rect 690 315 693 323
rect 1322 313 1356 316
rect 1370 313 1380 316
rect 1596 313 1613 316
rect 1634 315 1637 323
rect 1882 316 1885 323
rect 1826 313 1844 316
rect 1868 313 1885 316
rect 1364 303 1389 306
rect 1404 303 1469 306
rect 2004 303 2021 306
rect 2276 303 2293 306
rect 2402 303 2420 306
rect 14 267 2722 273
rect 1348 233 1381 236
rect 1428 233 1453 236
rect 2188 233 2205 236
rect 2236 233 2245 236
rect 194 216 197 225
rect 570 216 573 225
rect 722 216 725 225
rect 892 223 901 226
rect 932 223 965 226
rect 1322 223 1340 226
rect 1364 223 1373 226
rect 1450 223 1460 226
rect 1516 223 1525 226
rect 1988 223 1996 226
rect 2042 223 2060 226
rect 2074 223 2084 226
rect 1370 216 1373 223
rect 180 213 197 216
rect 212 213 221 216
rect 356 213 381 216
rect 556 213 573 216
rect 588 213 597 216
rect 636 213 661 216
rect 708 213 725 216
rect 740 213 749 216
rect 788 213 813 216
rect 844 213 853 216
rect 860 213 869 216
rect 890 213 916 216
rect 954 213 972 216
rect 1004 213 1013 216
rect 1018 213 1028 216
rect 1082 213 1108 216
rect 1370 213 1388 216
rect 1476 213 1485 216
rect 1522 213 1556 216
rect 1594 213 1613 216
rect 1644 213 1653 216
rect 186 203 196 206
rect 562 203 572 206
rect 850 205 853 213
rect 866 205 869 213
rect 1002 203 1036 206
rect 1066 203 1084 206
rect 1188 203 1196 206
rect 1250 203 1268 206
rect 1316 203 1333 206
rect 1580 203 1589 206
rect 1378 193 1388 196
rect 1610 195 1613 213
rect 1738 206 1741 214
rect 1746 213 1764 216
rect 1844 213 1853 216
rect 1948 213 1965 216
rect 1986 213 1997 216
rect 2018 213 2036 216
rect 1626 203 1636 206
rect 1738 203 1772 206
rect 1818 203 1836 206
rect 1884 203 1940 206
rect 1962 205 1965 213
rect 1994 205 1997 213
rect 2020 203 2029 206
rect 2044 203 2053 206
rect 2074 203 2077 214
rect 2106 213 2116 216
rect 2122 213 2140 216
rect 2274 203 2277 214
rect 2300 213 2317 216
rect 2364 213 2373 216
rect 2466 206 2469 214
rect 2532 213 2549 216
rect 2570 213 2596 216
rect 2308 203 2324 206
rect 2362 203 2372 206
rect 2466 203 2484 206
rect 2490 203 2500 206
rect 2514 203 2524 206
rect 2538 203 2548 206
rect 2570 205 2573 213
rect 1780 193 1829 196
rect 1850 193 1868 196
rect 2330 193 2340 196
rect 38 167 2698 173
rect 66 143 76 146
rect 1282 136 1285 145
rect 84 133 92 136
rect 210 126 213 135
rect 226 133 236 136
rect 362 126 365 135
rect 378 133 388 136
rect 514 126 517 135
rect 530 133 540 136
rect 666 126 669 135
rect 682 133 692 136
rect 818 126 821 135
rect 834 126 837 135
rect 962 126 965 135
rect 1084 133 1092 136
rect 1282 133 1292 136
rect 1386 133 1396 136
rect 1426 133 1444 136
rect 1458 133 1476 136
rect 100 123 109 126
rect 148 123 173 126
rect 204 123 213 126
rect 220 123 237 126
rect 300 123 325 126
rect 356 123 365 126
rect 372 123 389 126
rect 452 123 477 126
rect 508 123 517 126
rect 524 123 541 126
rect 556 123 565 126
rect 604 123 629 126
rect 660 123 669 126
rect 676 123 693 126
rect 756 123 781 126
rect 812 123 821 126
rect 828 123 837 126
rect 900 123 925 126
rect 956 123 965 126
rect 994 123 1004 126
rect 1228 123 1253 126
rect 1356 124 1372 127
rect 1412 123 1437 126
rect 1452 123 1469 126
rect 1482 125 1485 136
rect 1514 133 1548 136
rect 1596 133 1613 136
rect 1642 126 1645 135
rect 1668 133 1685 136
rect 1756 133 1773 136
rect 1794 126 1797 135
rect 1948 133 2005 136
rect 2026 133 2108 136
rect 1516 123 1549 126
rect 1628 123 1645 126
rect 1716 123 1733 126
rect 1762 123 1797 126
rect 2114 125 2117 136
rect 2228 133 2237 136
rect 2204 124 2220 127
rect 2226 123 2236 126
rect 234 115 237 123
rect 386 115 389 123
rect 538 115 541 123
rect 690 115 693 123
rect 1354 113 1364 116
rect 1668 113 1677 116
rect 1682 113 1708 116
rect 1722 113 1732 116
rect 1954 113 2004 116
rect 2122 113 2188 116
rect 2202 113 2212 116
rect 1348 103 1365 106
rect 2196 103 2213 106
rect 2845 76 2849 372
rect -102 -171 -98 72
rect 14 67 2722 73
rect 38 42 2698 57
rect 38 38 1224 42
rect 1228 38 2698 42
rect 38 37 2698 38
rect 14 13 2722 33
rect -68 -156 1185 -16
rect 1223 -171 1227 -23
rect 1249 -150 2750 -10
rect 2845 -170 2849 72
rect -98 -175 199 -171
rect 203 -175 499 -171
rect 803 -175 1227 -171
rect 1403 -174 1699 -170
rect 1703 -174 1999 -170
rect 2003 -174 2299 -170
rect 2303 -174 2599 -170
rect 2603 -174 2849 -170
rect 1223 -190 1227 -175
rect -1095 -917 -816 -222
rect 3570 -917 3853 -278
rect -1096 -1186 -164 -917
rect 2890 -1180 3853 -917
rect 2890 -1191 3851 -1180
<< m2contact >>
rect -101 2771 -97 2775
rect 199 2771 203 2775
rect 499 2771 503 2775
rect 799 2771 803 2775
rect 1347 2771 1351 2775
rect 1699 2771 1703 2775
rect 1999 2771 2003 2775
rect 2299 2771 2303 2775
rect 2599 2771 2603 2775
rect 2844 2771 2848 2775
rect -101 2472 -97 2476
rect 2844 2472 2848 2476
rect -101 2172 -97 2176
rect 2844 2172 2848 2176
rect -101 1872 -97 1876
rect 2844 1872 2848 1876
rect 2844 1572 2848 1576
rect -102 1272 -98 1276
rect 2844 1272 2848 1276
rect -102 972 -98 976
rect -102 672 -98 676
rect 2845 673 2849 677
rect -102 372 -98 376
rect 2845 372 2849 376
rect -102 72 -98 76
rect 2845 72 2849 76
rect 1224 38 1228 42
rect 1223 -23 1227 -19
rect -102 -175 -98 -171
rect 199 -175 203 -171
rect 499 -175 503 -171
rect 799 -175 803 -171
rect 1399 -174 1403 -170
rect 1699 -174 1703 -170
rect 1999 -174 2003 -170
rect 2299 -174 2303 -170
rect 2599 -174 2603 -170
<< metal2 >>
rect -100 2775 -97 2784
rect -109 2771 -101 2774
rect 134 2664 137 2783
rect 199 2775 202 2784
rect 435 2746 438 2783
rect 499 2775 502 2784
rect 735 2744 738 2784
rect 799 2775 802 2783
rect 1035 2746 1038 2783
rect 1112 2747 1115 2784
rect 1348 2775 1351 2783
rect 1700 2775 1703 2784
rect 1935 2736 1938 2785
rect 1999 2775 2002 2784
rect -26 2661 137 2664
rect 439 2733 1938 2736
rect -109 2537 -38 2540
rect -109 2472 -101 2475
rect -109 2236 -32 2239
rect -109 2172 -101 2175
rect -35 2097 -32 2236
rect -26 2137 -23 2661
rect -17 2186 -14 2651
rect -7 2207 -4 2643
rect 439 2638 442 2733
rect 2236 2727 2239 2785
rect 2299 2775 2302 2784
rect 474 2724 2239 2727
rect 474 2640 477 2724
rect 2535 2711 2538 2785
rect 2599 2775 2602 2783
rect 0 2635 442 2638
rect 458 2637 477 2640
rect 770 2708 2538 2711
rect 0 2407 3 2635
rect -17 2183 -8 2186
rect -26 2134 0 2137
rect -35 2094 3 2097
rect -109 1936 -9 1939
rect -110 1872 -101 1875
rect -109 1637 -23 1640
rect -108 1272 -102 1275
rect -26 1274 -23 1637
rect -109 1251 -18 1254
rect -21 1132 -18 1251
rect -12 1147 -9 1936
rect 0 1327 3 2094
rect -21 1129 -6 1132
rect -9 993 -6 1129
rect 1 1007 4 1268
rect -9 990 3 993
rect -108 972 -102 975
rect -109 950 -5 953
rect -8 808 -5 950
rect 0 817 3 990
rect -8 805 3 808
rect 0 737 3 805
rect -88 712 0 715
rect -108 672 -102 675
rect -88 653 -85 712
rect -110 650 -85 653
rect -108 372 -102 375
rect -88 353 -85 637
rect -110 350 -85 353
rect -80 532 0 535
rect -109 72 -102 75
rect -88 53 -85 335
rect -109 50 -85 53
rect -101 -184 -98 -175
rect -80 -185 -77 532
rect -74 332 0 335
rect -74 -159 -71 332
rect -68 173 0 176
rect -68 -153 -65 173
rect 14 13 34 2627
rect 38 37 58 2603
rect 66 2393 69 2406
rect 82 2403 85 2416
rect 82 2346 85 2366
rect 66 2333 69 2346
rect 74 2343 85 2346
rect 74 2296 77 2343
rect 82 2323 85 2336
rect 98 2333 101 2426
rect 178 2423 181 2546
rect 274 2533 277 2546
rect 226 2513 229 2526
rect 258 2476 261 2526
rect 250 2473 261 2476
rect 146 2393 149 2416
rect 186 2373 189 2416
rect 194 2406 197 2426
rect 194 2403 201 2406
rect 146 2323 149 2346
rect 162 2336 165 2356
rect 162 2333 173 2336
rect 74 2293 85 2296
rect 82 2236 85 2293
rect 170 2286 173 2333
rect 74 2233 85 2236
rect 162 2283 173 2286
rect 74 2213 77 2233
rect 106 2213 109 2226
rect 66 2183 69 2206
rect 66 2113 69 2136
rect 90 2133 93 2206
rect 114 2173 117 2216
rect 162 2186 165 2283
rect 186 2263 189 2326
rect 198 2306 201 2403
rect 210 2323 213 2426
rect 218 2393 221 2406
rect 226 2346 229 2416
rect 234 2353 237 2406
rect 218 2333 221 2346
rect 226 2343 245 2346
rect 226 2323 229 2343
rect 198 2303 205 2306
rect 202 2246 205 2303
rect 194 2243 205 2246
rect 170 2193 173 2216
rect 194 2203 197 2243
rect 218 2213 221 2226
rect 234 2223 237 2336
rect 242 2333 245 2343
rect 250 2273 253 2473
rect 266 2413 269 2426
rect 274 2403 277 2516
rect 282 2413 309 2416
rect 282 2403 293 2406
rect 290 2386 293 2403
rect 286 2383 293 2386
rect 258 2243 261 2336
rect 274 2256 277 2336
rect 286 2326 289 2383
rect 298 2333 301 2406
rect 306 2376 309 2413
rect 314 2403 317 2526
rect 306 2373 317 2376
rect 286 2323 293 2326
rect 270 2253 277 2256
rect 234 2213 245 2216
rect 162 2183 173 2186
rect 74 1743 77 2016
rect 138 2013 141 2126
rect 162 2116 165 2176
rect 170 2126 173 2183
rect 178 2133 181 2146
rect 210 2143 213 2206
rect 226 2193 229 2206
rect 234 2186 237 2213
rect 226 2183 237 2186
rect 170 2123 189 2126
rect 194 2123 197 2136
rect 162 2113 181 2116
rect 178 2036 181 2113
rect 178 2033 189 2036
rect 162 1973 165 2006
rect 186 1976 189 2033
rect 210 2013 213 2126
rect 226 2113 229 2183
rect 234 2123 237 2136
rect 242 2123 245 2206
rect 258 2193 261 2206
rect 250 2133 253 2176
rect 258 2133 261 2186
rect 270 2156 273 2253
rect 282 2213 285 2236
rect 266 2153 273 2156
rect 282 2153 285 2206
rect 250 2106 253 2126
rect 234 2013 237 2106
rect 246 2103 253 2106
rect 246 2026 249 2103
rect 246 2023 253 2026
rect 210 1983 213 2006
rect 178 1973 189 1976
rect 90 1896 93 1926
rect 122 1923 125 1936
rect 130 1923 133 1936
rect 90 1893 101 1896
rect 98 1826 101 1893
rect 90 1823 101 1826
rect 154 1823 157 1836
rect 90 1803 93 1823
rect 162 1816 165 1936
rect 130 1813 149 1816
rect 154 1813 165 1816
rect 90 1743 109 1746
rect 98 1613 101 1736
rect 106 1733 109 1743
rect 122 1703 125 1726
rect 130 1606 133 1636
rect 138 1623 141 1796
rect 146 1696 149 1806
rect 154 1793 157 1813
rect 170 1776 173 1926
rect 178 1843 181 1973
rect 186 1923 189 1946
rect 210 1933 213 1976
rect 226 1943 229 2006
rect 242 1993 245 2006
rect 226 1933 237 1936
rect 186 1823 205 1826
rect 194 1796 197 1816
rect 202 1803 205 1823
rect 186 1793 197 1796
rect 170 1773 181 1776
rect 162 1733 165 1746
rect 178 1743 181 1773
rect 154 1713 157 1726
rect 146 1693 153 1696
rect 150 1616 153 1693
rect 170 1666 173 1736
rect 186 1733 189 1793
rect 210 1756 213 1836
rect 178 1713 181 1726
rect 194 1716 197 1756
rect 202 1753 213 1756
rect 218 1753 221 1846
rect 202 1726 205 1753
rect 210 1733 213 1746
rect 202 1723 213 1726
rect 218 1723 221 1736
rect 226 1723 229 1926
rect 234 1836 237 1926
rect 242 1863 245 1956
rect 250 1923 253 2023
rect 258 1946 261 2126
rect 266 2123 269 2153
rect 274 2056 277 2136
rect 282 2113 285 2126
rect 290 2103 293 2323
rect 298 2066 301 2246
rect 306 2196 309 2366
rect 314 2323 317 2373
rect 322 2346 325 2426
rect 354 2413 357 2526
rect 370 2426 373 2546
rect 394 2476 397 2526
rect 450 2476 453 2536
rect 458 2533 461 2637
rect 482 2533 485 2546
rect 366 2423 373 2426
rect 386 2473 397 2476
rect 442 2473 453 2476
rect 466 2473 469 2526
rect 506 2506 509 2526
rect 506 2503 517 2506
rect 354 2363 357 2406
rect 366 2376 369 2423
rect 378 2403 381 2416
rect 386 2403 389 2473
rect 442 2426 445 2473
rect 474 2466 477 2496
rect 394 2413 397 2426
rect 434 2423 445 2426
rect 466 2463 477 2466
rect 366 2373 373 2376
rect 322 2343 333 2346
rect 314 2213 317 2226
rect 322 2213 325 2336
rect 330 2323 333 2343
rect 338 2333 341 2346
rect 338 2213 341 2286
rect 346 2243 349 2326
rect 354 2286 357 2336
rect 370 2333 373 2373
rect 394 2323 397 2346
rect 354 2283 365 2286
rect 362 2213 365 2283
rect 378 2216 381 2226
rect 370 2213 381 2216
rect 306 2193 313 2196
rect 310 2106 313 2193
rect 306 2103 313 2106
rect 306 2083 309 2103
rect 298 2063 309 2066
rect 274 2053 301 2056
rect 266 1966 269 1986
rect 274 1973 277 2046
rect 298 2013 301 2053
rect 266 1963 285 1966
rect 258 1943 277 1946
rect 258 1923 261 1943
rect 234 1833 245 1836
rect 242 1813 245 1833
rect 258 1813 261 1896
rect 266 1846 269 1936
rect 274 1933 277 1943
rect 274 1903 277 1926
rect 282 1913 285 1963
rect 306 1936 309 2063
rect 322 2056 325 2126
rect 318 2053 325 2056
rect 318 1966 321 2053
rect 338 1993 341 2186
rect 346 2143 349 2206
rect 370 2166 373 2206
rect 370 2163 389 2166
rect 354 2016 357 2106
rect 362 2043 365 2136
rect 386 2123 389 2163
rect 346 2013 357 2016
rect 370 2013 373 2086
rect 386 2013 389 2116
rect 394 2066 397 2176
rect 402 2086 405 2406
rect 410 2133 413 2206
rect 418 2183 421 2206
rect 402 2083 413 2086
rect 394 2063 401 2066
rect 346 1966 349 2013
rect 398 2006 401 2063
rect 410 2016 413 2083
rect 426 2033 429 2276
rect 434 2163 437 2423
rect 442 2276 445 2406
rect 450 2403 453 2416
rect 466 2406 469 2463
rect 474 2413 477 2426
rect 466 2403 477 2406
rect 450 2283 453 2326
rect 442 2273 453 2276
rect 442 2156 445 2216
rect 450 2173 453 2273
rect 458 2166 461 2336
rect 466 2313 469 2336
rect 474 2333 477 2346
rect 482 2323 485 2416
rect 490 2303 493 2476
rect 514 2446 517 2503
rect 498 2403 501 2446
rect 506 2443 517 2446
rect 506 2403 509 2443
rect 514 2413 517 2426
rect 546 2393 549 2406
rect 554 2366 557 2486
rect 562 2413 565 2576
rect 578 2533 581 2556
rect 626 2523 629 2546
rect 682 2533 685 2546
rect 666 2513 669 2526
rect 682 2493 685 2516
rect 714 2443 717 2546
rect 722 2503 725 2526
rect 730 2523 733 2536
rect 578 2413 589 2416
rect 562 2383 565 2406
rect 554 2363 561 2366
rect 466 2193 469 2216
rect 434 2153 445 2156
rect 410 2013 421 2016
rect 318 1963 325 1966
rect 290 1933 309 1936
rect 314 1933 317 1946
rect 290 1893 293 1933
rect 298 1913 301 1926
rect 306 1923 317 1926
rect 306 1903 309 1923
rect 322 1906 325 1963
rect 330 1963 349 1966
rect 354 2003 365 2006
rect 330 1933 333 1963
rect 330 1913 333 1926
rect 338 1906 341 1936
rect 314 1903 325 1906
rect 330 1903 341 1906
rect 266 1843 293 1846
rect 282 1823 285 1836
rect 274 1813 285 1816
rect 290 1806 293 1843
rect 298 1823 301 1846
rect 274 1803 293 1806
rect 298 1793 301 1806
rect 186 1713 197 1716
rect 210 1713 213 1723
rect 170 1663 181 1666
rect 106 1603 133 1606
rect 146 1613 153 1616
rect 162 1613 165 1626
rect 178 1616 181 1663
rect 186 1633 189 1713
rect 194 1623 197 1636
rect 178 1613 205 1616
rect 146 1593 149 1613
rect 210 1603 213 1646
rect 242 1643 245 1786
rect 226 1623 237 1626
rect 226 1613 229 1623
rect 242 1613 245 1636
rect 250 1623 253 1636
rect 258 1596 261 1786
rect 266 1603 269 1626
rect 274 1623 277 1736
rect 298 1733 301 1746
rect 282 1613 285 1636
rect 290 1633 293 1726
rect 306 1723 309 1816
rect 314 1733 317 1903
rect 330 1833 333 1903
rect 346 1896 349 1956
rect 338 1893 349 1896
rect 338 1813 341 1893
rect 346 1823 349 1886
rect 322 1743 333 1746
rect 298 1623 301 1636
rect 330 1633 333 1726
rect 314 1623 325 1626
rect 322 1606 325 1616
rect 306 1603 325 1606
rect 226 1593 237 1596
rect 258 1593 269 1596
rect 306 1593 309 1603
rect 82 1533 85 1546
rect 106 1476 109 1526
rect 162 1503 165 1526
rect 98 1473 109 1476
rect 98 1323 101 1473
rect 178 1436 181 1546
rect 130 1423 133 1436
rect 106 1146 109 1346
rect 130 1336 133 1416
rect 138 1406 141 1436
rect 146 1413 149 1426
rect 154 1413 157 1436
rect 178 1433 189 1436
rect 138 1403 157 1406
rect 154 1393 157 1403
rect 130 1333 149 1336
rect 154 1333 157 1346
rect 114 1213 117 1226
rect 106 1143 117 1146
rect 66 1013 69 1126
rect 82 1123 85 1136
rect 114 1096 117 1143
rect 130 1123 133 1326
rect 138 1316 141 1326
rect 146 1323 149 1333
rect 154 1316 157 1326
rect 138 1313 157 1316
rect 138 1223 141 1313
rect 146 1216 149 1226
rect 138 1213 149 1216
rect 154 1213 157 1226
rect 162 1213 165 1416
rect 178 1413 181 1426
rect 170 1283 173 1396
rect 162 1193 165 1206
rect 170 1136 173 1236
rect 178 1206 181 1306
rect 186 1233 189 1433
rect 202 1403 205 1526
rect 258 1513 261 1526
rect 266 1513 269 1593
rect 330 1583 333 1626
rect 338 1613 341 1806
rect 346 1573 349 1736
rect 354 1623 357 2003
rect 370 1956 373 1996
rect 378 1963 381 2006
rect 394 2003 401 2006
rect 370 1953 381 1956
rect 394 1953 397 2003
rect 362 1923 365 1936
rect 378 1933 381 1953
rect 362 1883 365 1916
rect 362 1833 365 1866
rect 362 1796 365 1816
rect 370 1813 373 1906
rect 378 1846 381 1926
rect 402 1923 405 1966
rect 378 1843 389 1846
rect 378 1823 381 1836
rect 362 1793 369 1796
rect 366 1736 369 1793
rect 362 1733 369 1736
rect 378 1733 381 1756
rect 362 1703 365 1733
rect 386 1723 389 1843
rect 394 1716 397 1826
rect 402 1793 405 1916
rect 410 1783 413 1996
rect 418 1813 421 2013
rect 426 1886 429 2006
rect 434 2003 437 2153
rect 450 2146 453 2166
rect 458 2163 469 2166
rect 442 2143 453 2146
rect 442 2003 445 2143
rect 426 1883 437 1886
rect 434 1753 437 1883
rect 442 1823 445 1996
rect 450 1983 453 2136
rect 458 1976 461 2156
rect 466 2146 469 2163
rect 466 2143 473 2146
rect 470 2036 473 2143
rect 482 2136 485 2216
rect 490 2183 493 2206
rect 498 2196 501 2356
rect 506 2323 509 2336
rect 522 2333 525 2356
rect 546 2323 549 2346
rect 558 2316 561 2363
rect 554 2313 561 2316
rect 514 2213 517 2306
rect 530 2213 533 2226
rect 498 2193 509 2196
rect 482 2133 493 2136
rect 466 2033 473 2036
rect 466 2013 469 2033
rect 482 2013 485 2126
rect 490 2083 493 2133
rect 506 2096 509 2193
rect 522 2133 525 2206
rect 554 2146 557 2313
rect 570 2156 573 2326
rect 586 2213 589 2386
rect 594 2323 605 2326
rect 610 2323 613 2406
rect 626 2403 629 2426
rect 634 2403 637 2416
rect 618 2306 621 2396
rect 626 2376 629 2396
rect 642 2393 645 2416
rect 658 2413 677 2416
rect 682 2413 685 2426
rect 626 2373 633 2376
rect 610 2303 621 2306
rect 610 2213 613 2303
rect 630 2296 633 2373
rect 642 2343 645 2386
rect 650 2336 653 2376
rect 626 2293 633 2296
rect 642 2333 653 2336
rect 626 2243 629 2293
rect 626 2226 629 2236
rect 618 2223 629 2226
rect 618 2213 621 2223
rect 634 2213 637 2226
rect 578 2193 581 2206
rect 570 2153 581 2156
rect 554 2143 573 2146
rect 498 2093 509 2096
rect 498 2076 501 2093
rect 490 2073 501 2076
rect 450 1973 461 1976
rect 450 1863 453 1973
rect 458 1843 461 1966
rect 466 1836 469 2006
rect 474 2003 485 2006
rect 490 1973 493 2073
rect 538 2066 541 2136
rect 562 2123 565 2136
rect 570 2073 573 2143
rect 578 2106 581 2153
rect 586 2123 589 2206
rect 578 2103 585 2106
rect 514 2063 541 2066
rect 474 1886 477 1926
rect 482 1913 485 1926
rect 474 1883 485 1886
rect 442 1763 445 1806
rect 378 1713 397 1716
rect 378 1656 381 1713
rect 370 1653 381 1656
rect 362 1613 365 1626
rect 354 1593 357 1606
rect 370 1596 373 1653
rect 378 1613 381 1626
rect 386 1603 389 1636
rect 394 1603 397 1616
rect 402 1603 405 1616
rect 370 1593 389 1596
rect 282 1523 293 1526
rect 274 1486 277 1506
rect 266 1483 277 1486
rect 266 1466 269 1483
rect 258 1463 269 1466
rect 258 1403 261 1463
rect 282 1446 285 1516
rect 274 1443 285 1446
rect 210 1303 213 1326
rect 218 1313 221 1396
rect 266 1323 269 1406
rect 274 1323 277 1443
rect 290 1356 293 1523
rect 306 1523 333 1526
rect 298 1436 301 1516
rect 306 1513 309 1523
rect 314 1486 317 1506
rect 322 1503 325 1516
rect 330 1513 333 1523
rect 330 1486 333 1506
rect 314 1483 333 1486
rect 298 1433 309 1436
rect 282 1353 293 1356
rect 282 1293 285 1353
rect 290 1343 301 1346
rect 186 1213 189 1226
rect 178 1203 189 1206
rect 162 1133 173 1136
rect 162 1123 165 1133
rect 106 1093 117 1096
rect 66 993 69 1006
rect 66 976 69 986
rect 74 983 77 1016
rect 106 1013 109 1093
rect 122 1043 149 1046
rect 122 1003 125 1043
rect 146 1026 149 1043
rect 130 1013 133 1026
rect 146 1023 157 1026
rect 130 993 133 1006
rect 66 973 85 976
rect 82 923 85 973
rect 106 923 109 986
rect 138 966 141 1016
rect 146 993 149 1016
rect 154 996 157 1023
rect 162 1003 165 1086
rect 170 1076 173 1126
rect 178 1083 181 1126
rect 186 1123 189 1196
rect 202 1176 205 1206
rect 198 1173 205 1176
rect 198 1086 201 1173
rect 226 1126 229 1216
rect 266 1133 269 1196
rect 282 1153 285 1286
rect 290 1203 293 1336
rect 298 1306 301 1336
rect 306 1333 309 1433
rect 338 1336 341 1526
rect 354 1513 357 1586
rect 362 1533 365 1546
rect 386 1533 389 1593
rect 362 1456 365 1526
rect 354 1453 365 1456
rect 314 1333 325 1336
rect 330 1333 341 1336
rect 346 1333 349 1346
rect 314 1313 317 1326
rect 298 1303 317 1306
rect 298 1213 301 1296
rect 330 1223 333 1333
rect 322 1193 325 1216
rect 218 1123 229 1126
rect 198 1083 205 1086
rect 170 1073 181 1076
rect 170 1003 173 1016
rect 178 1003 181 1073
rect 202 1026 205 1083
rect 186 1013 189 1026
rect 194 1023 205 1026
rect 154 993 165 996
rect 138 963 149 966
rect 146 933 149 963
rect 122 913 125 926
rect 74 813 85 816
rect 130 793 133 816
rect 74 663 77 726
rect 130 723 133 746
rect 74 613 85 616
rect 82 573 85 613
rect 130 603 133 616
rect 154 576 157 926
rect 162 923 165 993
rect 194 973 197 1023
rect 202 993 205 1016
rect 210 993 213 1006
rect 218 1003 221 1123
rect 242 1076 245 1126
rect 290 1123 293 1136
rect 314 1123 317 1156
rect 242 1073 253 1076
rect 226 996 229 1006
rect 234 1003 237 1016
rect 242 1013 245 1036
rect 242 996 245 1006
rect 250 1003 253 1073
rect 258 1013 261 1046
rect 226 993 245 996
rect 170 913 173 926
rect 226 913 229 926
rect 250 876 253 976
rect 266 953 269 1006
rect 274 946 277 1036
rect 282 1013 285 1106
rect 322 1103 325 1186
rect 290 1013 293 1046
rect 298 966 301 1026
rect 306 1023 325 1026
rect 306 1003 309 1016
rect 314 1003 317 1016
rect 298 963 309 966
rect 266 943 277 946
rect 266 933 269 943
rect 274 923 277 936
rect 290 913 293 926
rect 298 913 301 956
rect 234 873 253 876
rect 186 816 189 836
rect 170 803 173 816
rect 178 813 189 816
rect 170 713 173 736
rect 178 726 181 813
rect 186 793 189 806
rect 186 733 189 746
rect 194 733 197 756
rect 210 733 213 816
rect 178 723 189 726
rect 186 656 189 723
rect 178 576 181 656
rect 186 653 213 656
rect 138 573 157 576
rect 170 573 181 576
rect 66 496 69 536
rect 90 513 93 526
rect 138 496 141 573
rect 146 523 149 546
rect 170 533 173 573
rect 186 533 189 576
rect 202 533 205 606
rect 210 526 213 653
rect 218 536 221 826
rect 234 653 237 873
rect 306 826 309 963
rect 314 933 317 996
rect 322 913 325 1016
rect 330 913 333 1216
rect 346 1193 349 1206
rect 354 1183 357 1453
rect 378 1423 381 1526
rect 362 1313 365 1326
rect 370 1296 373 1336
rect 366 1293 373 1296
rect 366 1226 369 1293
rect 366 1223 373 1226
rect 370 1203 373 1223
rect 378 1196 381 1416
rect 386 1306 389 1526
rect 394 1413 397 1586
rect 410 1566 413 1726
rect 442 1723 445 1746
rect 418 1593 421 1616
rect 426 1603 429 1646
rect 402 1563 413 1566
rect 402 1496 405 1563
rect 410 1503 413 1556
rect 426 1523 429 1546
rect 434 1523 437 1706
rect 402 1493 413 1496
rect 410 1436 413 1493
rect 410 1433 417 1436
rect 394 1323 397 1406
rect 386 1303 393 1306
rect 338 973 341 1146
rect 338 933 341 956
rect 346 916 349 1086
rect 354 1023 357 1176
rect 338 913 349 916
rect 354 926 357 1016
rect 362 936 365 1196
rect 370 1193 381 1196
rect 370 1153 373 1193
rect 378 1133 381 1166
rect 390 1146 393 1303
rect 386 1143 393 1146
rect 402 1143 405 1426
rect 414 1386 417 1433
rect 410 1383 417 1386
rect 410 1333 413 1383
rect 426 1353 429 1416
rect 442 1403 445 1716
rect 450 1576 453 1836
rect 458 1833 469 1836
rect 458 1743 461 1833
rect 466 1733 469 1826
rect 474 1786 477 1866
rect 482 1813 485 1883
rect 490 1803 493 1926
rect 498 1896 501 2006
rect 514 1993 517 2063
rect 562 2036 565 2056
rect 554 2033 565 2036
rect 538 2003 541 2016
rect 506 1933 509 1976
rect 514 1943 517 1986
rect 554 1966 557 2033
rect 582 2016 585 2103
rect 578 2013 585 2016
rect 578 1993 581 2013
rect 554 1963 565 1966
rect 530 1943 557 1946
rect 498 1893 509 1896
rect 506 1846 509 1893
rect 498 1843 509 1846
rect 498 1793 501 1843
rect 474 1783 501 1786
rect 482 1733 485 1756
rect 458 1723 477 1726
rect 474 1706 477 1716
rect 482 1713 485 1726
rect 490 1713 493 1766
rect 498 1723 501 1783
rect 506 1716 509 1826
rect 522 1816 525 1936
rect 530 1896 533 1943
rect 538 1906 541 1936
rect 546 1923 549 1936
rect 554 1913 557 1926
rect 538 1903 549 1906
rect 530 1893 541 1896
rect 538 1823 541 1893
rect 546 1836 549 1903
rect 562 1873 565 1963
rect 570 1933 573 1956
rect 586 1936 589 1966
rect 594 1943 597 2016
rect 578 1926 581 1936
rect 586 1933 597 1936
rect 602 1933 605 2196
rect 610 1973 613 2156
rect 610 1933 613 1946
rect 570 1923 581 1926
rect 586 1913 589 1926
rect 594 1923 605 1926
rect 610 1913 613 1926
rect 618 1923 621 2176
rect 626 2113 629 2166
rect 642 2153 645 2333
rect 666 2306 669 2396
rect 674 2346 677 2406
rect 682 2393 685 2406
rect 698 2356 701 2426
rect 706 2366 709 2426
rect 714 2423 717 2436
rect 730 2413 733 2516
rect 746 2506 749 2526
rect 742 2503 749 2506
rect 742 2436 745 2503
rect 754 2466 757 2536
rect 770 2533 773 2708
rect 2834 2698 2837 2785
rect 2848 2772 2858 2775
rect 850 2695 2837 2698
rect 802 2533 805 2556
rect 818 2533 821 2576
rect 850 2553 853 2695
rect 930 2683 2788 2686
rect 930 2640 933 2683
rect 978 2670 2777 2673
rect 978 2640 981 2670
rect 930 2637 949 2640
rect 842 2533 845 2546
rect 858 2533 861 2566
rect 922 2546 925 2566
rect 762 2476 765 2526
rect 762 2473 773 2476
rect 754 2463 765 2466
rect 742 2433 749 2436
rect 746 2413 749 2433
rect 714 2373 717 2406
rect 706 2363 717 2366
rect 698 2353 709 2356
rect 674 2343 701 2346
rect 658 2303 669 2306
rect 682 2333 701 2336
rect 658 2213 661 2303
rect 666 2213 669 2236
rect 674 2213 677 2226
rect 658 2153 661 2206
rect 674 2133 677 2166
rect 642 2123 653 2126
rect 650 2093 653 2123
rect 626 1896 629 2046
rect 650 2036 653 2076
rect 634 1943 637 2036
rect 650 2033 661 2036
rect 674 2033 677 2116
rect 682 2113 685 2333
rect 698 2253 701 2326
rect 706 2323 709 2353
rect 714 2313 717 2363
rect 738 2333 741 2406
rect 754 2393 757 2426
rect 762 2413 765 2463
rect 762 2386 765 2406
rect 754 2383 765 2386
rect 754 2346 757 2383
rect 770 2363 773 2473
rect 826 2453 829 2526
rect 842 2443 845 2516
rect 858 2486 861 2526
rect 882 2523 885 2546
rect 922 2543 929 2546
rect 858 2483 869 2486
rect 778 2403 781 2426
rect 786 2413 789 2426
rect 802 2413 805 2426
rect 834 2413 837 2426
rect 746 2343 757 2346
rect 746 2293 749 2343
rect 754 2333 797 2336
rect 762 2303 765 2316
rect 770 2303 773 2316
rect 786 2303 789 2316
rect 762 2266 765 2286
rect 754 2263 765 2266
rect 690 2113 693 2156
rect 698 2133 701 2246
rect 706 2223 725 2226
rect 682 2093 685 2106
rect 618 1893 629 1896
rect 546 1833 557 1836
rect 546 1816 549 1826
rect 522 1813 533 1816
rect 538 1813 549 1816
rect 514 1803 525 1806
rect 514 1733 517 1746
rect 498 1713 509 1716
rect 498 1706 501 1713
rect 466 1576 469 1706
rect 474 1703 501 1706
rect 474 1603 477 1626
rect 450 1573 461 1576
rect 466 1573 477 1576
rect 458 1553 461 1573
rect 474 1533 477 1573
rect 482 1553 485 1656
rect 522 1613 525 1786
rect 530 1736 533 1813
rect 546 1763 549 1813
rect 554 1803 557 1833
rect 618 1826 621 1893
rect 634 1826 637 1936
rect 642 1913 645 2026
rect 658 1986 661 2033
rect 674 2013 685 2016
rect 690 2006 693 2026
rect 698 2013 701 2126
rect 706 2113 709 2223
rect 722 2216 725 2223
rect 722 2213 733 2216
rect 730 2193 733 2213
rect 714 2133 717 2176
rect 754 2166 757 2263
rect 770 2193 773 2206
rect 754 2163 765 2166
rect 714 2113 717 2126
rect 738 2023 741 2126
rect 762 2076 765 2163
rect 754 2073 765 2076
rect 690 2003 701 2006
rect 650 1983 661 1986
rect 650 1906 653 1983
rect 658 1913 661 1936
rect 666 1933 669 1966
rect 682 1933 685 1996
rect 698 1943 701 1956
rect 682 1906 685 1926
rect 650 1903 661 1906
rect 618 1823 629 1826
rect 634 1823 653 1826
rect 570 1813 581 1816
rect 602 1793 605 1806
rect 578 1743 581 1756
rect 586 1743 589 1776
rect 530 1733 549 1736
rect 546 1726 549 1733
rect 538 1606 541 1726
rect 546 1723 557 1726
rect 562 1693 565 1736
rect 594 1666 597 1756
rect 602 1703 605 1786
rect 610 1733 613 1806
rect 626 1783 629 1823
rect 618 1733 629 1736
rect 610 1713 613 1726
rect 618 1716 621 1726
rect 634 1723 637 1806
rect 642 1733 645 1806
rect 650 1803 653 1823
rect 618 1713 637 1716
rect 626 1683 629 1713
rect 586 1663 597 1666
rect 490 1533 493 1606
rect 538 1603 549 1606
rect 554 1603 557 1636
rect 538 1556 541 1596
rect 546 1563 549 1603
rect 570 1593 573 1616
rect 538 1553 549 1556
rect 578 1553 581 1616
rect 586 1583 589 1663
rect 602 1613 605 1646
rect 634 1576 637 1706
rect 642 1603 645 1636
rect 650 1583 653 1766
rect 658 1753 661 1903
rect 674 1903 685 1906
rect 674 1836 677 1903
rect 674 1833 685 1836
rect 666 1813 677 1816
rect 666 1783 669 1796
rect 658 1703 661 1716
rect 666 1703 669 1716
rect 674 1713 677 1806
rect 682 1773 685 1833
rect 690 1783 693 1936
rect 706 1923 709 1976
rect 754 1973 757 2073
rect 770 2066 773 2136
rect 778 2123 781 2276
rect 786 2213 789 2296
rect 794 2213 797 2333
rect 802 2273 805 2366
rect 834 2326 837 2406
rect 842 2383 845 2406
rect 866 2383 869 2483
rect 810 2323 837 2326
rect 794 2196 797 2206
rect 802 2203 805 2236
rect 810 2213 813 2266
rect 826 2233 829 2316
rect 834 2303 837 2316
rect 842 2283 845 2366
rect 842 2233 845 2256
rect 826 2223 845 2226
rect 826 2213 829 2223
rect 794 2193 821 2196
rect 714 1933 717 1966
rect 762 1963 765 2066
rect 770 2063 781 2066
rect 786 2063 789 2186
rect 834 2116 837 2136
rect 770 2003 773 2016
rect 778 2003 781 2063
rect 786 2013 789 2026
rect 794 2003 797 2086
rect 810 2023 813 2116
rect 826 2113 837 2116
rect 826 2066 829 2113
rect 826 2063 837 2066
rect 834 2013 837 2063
rect 762 1933 765 1956
rect 706 1833 725 1836
rect 706 1813 709 1833
rect 698 1793 701 1806
rect 706 1783 709 1806
rect 682 1653 685 1736
rect 690 1703 693 1726
rect 698 1593 701 1606
rect 706 1583 709 1686
rect 538 1496 541 1546
rect 546 1533 549 1553
rect 546 1513 549 1526
rect 562 1506 565 1526
rect 530 1493 541 1496
rect 546 1503 565 1506
rect 450 1393 453 1406
rect 386 1126 389 1143
rect 402 1126 405 1136
rect 370 1083 373 1126
rect 382 1123 389 1126
rect 394 1123 405 1126
rect 410 1123 413 1216
rect 418 1156 421 1206
rect 426 1173 429 1326
rect 434 1223 437 1236
rect 434 1193 437 1216
rect 418 1153 429 1156
rect 382 1076 385 1123
rect 418 1103 421 1136
rect 378 1073 385 1076
rect 370 943 373 1026
rect 378 1013 381 1073
rect 402 1013 405 1026
rect 426 1013 429 1153
rect 434 1113 437 1136
rect 442 1133 445 1306
rect 450 1183 453 1236
rect 458 1216 461 1336
rect 466 1303 469 1316
rect 474 1313 477 1326
rect 466 1223 469 1236
rect 458 1213 469 1216
rect 466 1203 469 1213
rect 474 1193 477 1306
rect 378 993 381 1006
rect 362 933 381 936
rect 354 923 373 926
rect 338 903 341 913
rect 346 883 349 906
rect 302 823 309 826
rect 282 803 285 816
rect 302 736 305 823
rect 258 716 261 736
rect 250 713 261 716
rect 250 636 253 713
rect 250 633 261 636
rect 226 593 229 616
rect 258 613 261 633
rect 266 603 269 726
rect 274 723 277 736
rect 302 733 309 736
rect 314 733 317 816
rect 322 763 325 836
rect 346 813 349 826
rect 306 716 309 733
rect 306 713 313 716
rect 274 556 277 626
rect 290 623 293 636
rect 298 613 301 706
rect 290 593 293 606
rect 310 576 313 713
rect 330 623 333 736
rect 346 733 349 806
rect 354 803 357 923
rect 362 893 365 916
rect 378 883 381 933
rect 386 856 389 926
rect 394 916 397 986
rect 402 933 405 956
rect 394 913 405 916
rect 394 893 397 906
rect 402 876 405 913
rect 370 853 389 856
rect 394 873 405 876
rect 362 813 365 826
rect 370 803 373 853
rect 354 703 357 736
rect 378 733 381 816
rect 386 813 389 826
rect 394 803 397 873
rect 402 803 405 816
rect 410 776 413 946
rect 418 813 421 976
rect 426 963 429 1006
rect 434 1003 437 1036
rect 442 983 445 1126
rect 450 1013 453 1156
rect 458 1113 461 1166
rect 466 1123 469 1136
rect 474 1016 477 1146
rect 482 1103 485 1356
rect 490 1263 493 1416
rect 530 1413 533 1493
rect 498 1356 501 1406
rect 530 1366 533 1386
rect 530 1363 537 1366
rect 498 1353 509 1356
rect 498 1303 501 1316
rect 506 1313 509 1353
rect 522 1323 525 1336
rect 514 1236 517 1306
rect 522 1303 525 1316
rect 534 1296 537 1363
rect 506 1233 517 1236
rect 530 1293 537 1296
rect 506 1206 509 1233
rect 514 1213 517 1226
rect 490 1163 493 1206
rect 506 1203 517 1206
rect 490 1133 493 1156
rect 498 1133 501 1146
rect 458 1013 477 1016
rect 490 1013 493 1126
rect 498 1113 501 1126
rect 506 1033 509 1186
rect 514 1123 517 1203
rect 522 1166 525 1216
rect 530 1173 533 1293
rect 538 1213 541 1236
rect 522 1163 533 1166
rect 522 1133 525 1156
rect 498 1013 501 1026
rect 450 993 453 1006
rect 458 976 461 1006
rect 466 983 469 1006
rect 442 973 461 976
rect 442 933 445 973
rect 474 956 477 996
rect 522 983 525 1116
rect 530 1076 533 1163
rect 538 1133 541 1146
rect 538 1113 541 1126
rect 530 1073 541 1076
rect 530 993 533 1006
rect 538 993 541 1073
rect 474 953 493 956
rect 426 793 429 896
rect 434 803 437 896
rect 410 773 421 776
rect 378 703 381 716
rect 394 623 397 726
rect 402 693 405 766
rect 418 636 421 773
rect 442 733 445 816
rect 458 806 461 926
rect 490 896 493 953
rect 514 933 517 946
rect 482 893 493 896
rect 482 826 485 893
rect 482 823 493 826
rect 458 803 469 806
rect 410 633 421 636
rect 354 593 357 616
rect 378 583 381 606
rect 394 593 397 606
rect 410 593 413 633
rect 418 603 421 616
rect 310 573 325 576
rect 266 553 277 556
rect 218 533 237 536
rect 202 523 213 526
rect 66 493 77 496
rect 138 493 157 496
rect 74 446 77 493
rect 66 443 77 446
rect 66 413 69 443
rect 130 393 133 416
rect 66 323 69 336
rect 130 323 133 346
rect 66 143 69 196
rect 74 173 77 216
rect 130 193 133 216
rect 106 123 109 146
rect 122 133 125 146
rect 154 143 157 493
rect 170 403 173 426
rect 186 416 189 426
rect 202 416 205 523
rect 186 413 205 416
rect 218 413 221 426
rect 186 393 189 406
rect 170 333 181 336
rect 186 333 189 346
rect 194 326 197 413
rect 186 323 197 326
rect 186 226 189 323
rect 218 316 221 406
rect 226 363 229 416
rect 234 393 237 533
rect 242 513 245 536
rect 266 336 269 553
rect 282 533 285 546
rect 282 513 285 526
rect 298 486 301 536
rect 322 513 325 573
rect 298 483 309 486
rect 282 393 285 416
rect 306 373 309 483
rect 322 386 325 406
rect 314 383 325 386
rect 210 313 221 316
rect 226 316 229 336
rect 258 323 261 336
rect 266 333 277 336
rect 226 313 237 316
rect 210 296 213 313
rect 202 293 213 296
rect 202 246 205 293
rect 202 243 213 246
rect 186 223 205 226
rect 170 173 173 206
rect 186 193 189 206
rect 202 196 205 223
rect 210 206 213 243
rect 218 213 221 306
rect 234 266 237 313
rect 226 263 237 266
rect 226 213 229 263
rect 210 203 221 206
rect 202 193 213 196
rect 170 123 173 146
rect 210 126 213 193
rect 218 163 221 203
rect 266 176 269 326
rect 274 293 277 333
rect 282 323 285 356
rect 298 326 301 336
rect 306 333 309 366
rect 290 323 301 326
rect 314 323 317 383
rect 330 353 333 416
rect 338 383 341 526
rect 346 423 349 436
rect 346 393 349 406
rect 354 403 357 426
rect 378 423 381 476
rect 394 423 397 526
rect 402 523 405 566
rect 426 563 429 606
rect 442 583 445 616
rect 450 446 453 796
rect 466 756 469 803
rect 458 753 469 756
rect 458 723 461 753
rect 482 736 485 806
rect 490 796 493 823
rect 498 803 501 836
rect 506 813 509 926
rect 522 823 525 956
rect 530 906 533 976
rect 538 933 541 946
rect 546 933 549 1503
rect 554 1403 557 1456
rect 562 1386 565 1416
rect 594 1413 597 1566
rect 602 1533 605 1576
rect 634 1573 661 1576
rect 602 1503 605 1526
rect 650 1523 653 1536
rect 658 1533 661 1573
rect 714 1563 717 1826
rect 722 1703 725 1826
rect 730 1693 733 1846
rect 738 1733 741 1926
rect 770 1916 773 1946
rect 766 1913 773 1916
rect 766 1846 769 1913
rect 766 1843 773 1846
rect 762 1813 765 1826
rect 746 1803 757 1806
rect 770 1803 773 1843
rect 778 1823 781 1976
rect 786 1913 789 1926
rect 778 1796 781 1816
rect 786 1803 789 1816
rect 770 1793 781 1796
rect 738 1633 741 1726
rect 746 1713 749 1726
rect 762 1703 765 1726
rect 770 1703 773 1793
rect 722 1603 725 1616
rect 738 1613 741 1626
rect 658 1483 661 1526
rect 682 1493 685 1526
rect 690 1513 693 1526
rect 558 1383 565 1386
rect 558 1246 561 1383
rect 570 1313 573 1406
rect 558 1243 565 1246
rect 554 1213 557 1226
rect 562 1213 565 1243
rect 562 1193 565 1206
rect 554 1063 557 1176
rect 570 1133 573 1306
rect 578 1303 597 1306
rect 578 1213 581 1303
rect 602 1213 605 1336
rect 626 1326 629 1416
rect 634 1403 637 1476
rect 690 1413 693 1426
rect 698 1406 701 1506
rect 706 1473 709 1546
rect 714 1466 717 1556
rect 722 1506 725 1576
rect 730 1523 733 1606
rect 754 1603 757 1636
rect 778 1613 781 1626
rect 738 1543 741 1566
rect 722 1503 729 1506
rect 642 1363 645 1406
rect 690 1403 701 1406
rect 706 1463 717 1466
rect 626 1323 637 1326
rect 690 1323 693 1403
rect 610 1296 613 1316
rect 610 1293 617 1296
rect 614 1226 617 1293
rect 634 1256 637 1323
rect 610 1223 617 1226
rect 626 1253 637 1256
rect 562 1096 565 1126
rect 570 1113 573 1126
rect 562 1093 573 1096
rect 562 1056 565 1093
rect 554 1053 565 1056
rect 554 1003 557 1053
rect 578 1043 581 1206
rect 586 1153 589 1206
rect 594 1163 597 1206
rect 586 1126 589 1146
rect 586 1123 593 1126
rect 590 1056 593 1123
rect 586 1053 593 1056
rect 586 1036 589 1053
rect 562 1013 565 1036
rect 570 1033 589 1036
rect 562 993 565 1006
rect 570 973 573 1033
rect 578 1023 589 1026
rect 594 953 597 1016
rect 602 1013 605 1206
rect 610 1113 613 1223
rect 618 1193 621 1206
rect 626 1203 629 1253
rect 698 1236 701 1396
rect 706 1333 709 1463
rect 726 1456 729 1503
rect 738 1486 741 1536
rect 746 1513 749 1576
rect 738 1483 749 1486
rect 722 1453 729 1456
rect 722 1426 725 1453
rect 718 1423 725 1426
rect 718 1316 721 1423
rect 714 1313 721 1316
rect 714 1256 717 1313
rect 730 1273 733 1416
rect 746 1413 749 1483
rect 754 1453 757 1586
rect 794 1563 797 1996
rect 810 1983 813 2006
rect 842 1976 845 2216
rect 850 2213 853 2306
rect 858 2303 861 2336
rect 866 2213 869 2316
rect 874 2286 877 2456
rect 882 2423 885 2496
rect 926 2486 929 2543
rect 946 2533 949 2637
rect 962 2637 981 2640
rect 1042 2661 2767 2664
rect 962 2533 965 2637
rect 986 2533 989 2566
rect 1042 2563 1045 2661
rect 1146 2653 2759 2656
rect 922 2483 929 2486
rect 882 2303 885 2416
rect 898 2413 901 2446
rect 906 2403 909 2456
rect 922 2403 925 2483
rect 938 2453 941 2526
rect 938 2333 941 2386
rect 874 2283 881 2286
rect 878 2206 881 2283
rect 890 2253 893 2316
rect 898 2303 901 2316
rect 906 2293 909 2326
rect 914 2313 925 2316
rect 930 2306 933 2326
rect 914 2303 933 2306
rect 930 2223 933 2236
rect 938 2216 941 2226
rect 874 2203 881 2206
rect 874 2146 877 2203
rect 874 2143 893 2146
rect 858 2056 861 2136
rect 890 2096 893 2143
rect 906 2123 909 2206
rect 930 2196 933 2216
rect 938 2213 949 2216
rect 954 2213 957 2526
rect 970 2443 973 2526
rect 1034 2523 1037 2546
rect 1074 2533 1077 2566
rect 1090 2533 1093 2576
rect 1114 2533 1117 2546
rect 1074 2523 1085 2526
rect 970 2393 973 2416
rect 1002 2383 1005 2416
rect 1010 2413 1013 2426
rect 970 2306 973 2326
rect 970 2303 981 2306
rect 978 2226 981 2303
rect 1010 2276 1013 2406
rect 1018 2376 1021 2446
rect 1034 2393 1037 2406
rect 1018 2373 1029 2376
rect 970 2223 981 2226
rect 1002 2273 1013 2276
rect 926 2193 933 2196
rect 926 2116 929 2193
rect 938 2123 941 2166
rect 946 2123 949 2213
rect 954 2203 965 2206
rect 970 2193 973 2223
rect 978 2193 981 2206
rect 1002 2203 1005 2273
rect 1026 2266 1029 2373
rect 1042 2333 1045 2406
rect 1018 2263 1029 2266
rect 1018 2216 1021 2263
rect 1042 2223 1045 2326
rect 1058 2313 1061 2496
rect 1098 2446 1101 2526
rect 1122 2523 1125 2536
rect 1146 2533 1149 2653
rect 1218 2645 2752 2648
rect 1218 2576 1221 2645
rect 1346 2637 2745 2640
rect 1210 2573 1221 2576
rect 1162 2533 1165 2556
rect 1194 2533 1197 2546
rect 1210 2533 1213 2573
rect 1138 2493 1141 2516
rect 1098 2443 1109 2446
rect 1074 2256 1077 2416
rect 1106 2396 1109 2443
rect 1122 2403 1125 2416
rect 1058 2253 1077 2256
rect 1098 2393 1109 2396
rect 1010 2193 1013 2216
rect 1018 2213 1029 2216
rect 954 2133 957 2166
rect 926 2113 933 2116
rect 850 2053 861 2056
rect 882 2093 893 2096
rect 850 1983 853 2053
rect 802 1916 805 1936
rect 810 1933 813 1966
rect 818 1923 821 1976
rect 842 1973 853 1976
rect 834 1933 837 1946
rect 842 1933 845 1956
rect 850 1926 853 1973
rect 842 1923 853 1926
rect 802 1913 809 1916
rect 806 1836 809 1913
rect 802 1833 809 1836
rect 802 1813 805 1833
rect 818 1773 821 1856
rect 834 1803 837 1816
rect 842 1786 845 1923
rect 858 1903 861 2006
rect 874 1933 877 1986
rect 882 1973 885 2093
rect 930 2046 933 2113
rect 930 2043 941 2046
rect 890 2003 893 2036
rect 906 1983 909 2006
rect 938 1996 941 2043
rect 922 1993 941 1996
rect 954 1993 957 2016
rect 898 1923 901 1946
rect 850 1796 853 1816
rect 850 1793 861 1796
rect 842 1783 853 1786
rect 802 1543 805 1616
rect 754 1413 757 1426
rect 754 1393 757 1406
rect 762 1333 765 1436
rect 770 1396 773 1416
rect 778 1403 781 1436
rect 786 1426 789 1526
rect 802 1483 805 1536
rect 786 1423 805 1426
rect 786 1396 789 1406
rect 770 1393 789 1396
rect 714 1253 725 1256
rect 650 1223 653 1236
rect 698 1233 717 1236
rect 618 1106 621 1186
rect 626 1146 629 1196
rect 634 1186 637 1206
rect 642 1193 645 1216
rect 650 1186 653 1216
rect 634 1183 653 1186
rect 634 1153 637 1183
rect 626 1143 637 1146
rect 614 1103 621 1106
rect 614 1026 617 1103
rect 626 1093 629 1106
rect 610 1023 617 1026
rect 602 946 605 1006
rect 610 963 613 1023
rect 626 1006 629 1046
rect 634 1033 637 1143
rect 642 1113 645 1166
rect 658 1156 661 1206
rect 706 1193 709 1206
rect 714 1193 717 1233
rect 722 1213 725 1253
rect 730 1206 733 1266
rect 738 1213 741 1326
rect 754 1246 757 1326
rect 770 1266 773 1326
rect 746 1243 757 1246
rect 762 1263 773 1266
rect 722 1203 733 1206
rect 690 1183 709 1186
rect 738 1183 741 1206
rect 746 1203 749 1243
rect 754 1213 757 1226
rect 762 1183 765 1263
rect 682 1156 685 1176
rect 658 1153 685 1156
rect 690 1153 693 1183
rect 738 1153 757 1156
rect 770 1153 773 1256
rect 778 1156 781 1366
rect 786 1253 789 1356
rect 794 1303 797 1416
rect 802 1293 805 1423
rect 802 1263 805 1286
rect 794 1213 797 1226
rect 802 1203 805 1246
rect 778 1153 789 1156
rect 650 1123 653 1136
rect 658 1093 661 1136
rect 666 1113 669 1126
rect 618 993 621 1006
rect 626 1003 637 1006
rect 626 953 629 996
rect 562 943 581 946
rect 562 933 565 943
rect 546 923 557 926
rect 530 903 541 906
rect 538 816 541 903
rect 562 833 565 926
rect 522 813 541 816
rect 562 813 565 826
rect 490 793 501 796
rect 466 683 469 736
rect 482 733 493 736
rect 474 703 477 726
rect 482 696 485 726
rect 474 693 485 696
rect 466 616 469 626
rect 458 613 469 616
rect 474 613 477 693
rect 458 573 461 613
rect 466 546 469 606
rect 482 583 485 686
rect 490 653 493 726
rect 498 723 501 793
rect 498 693 501 716
rect 506 686 509 736
rect 514 696 517 756
rect 522 733 525 813
rect 570 803 573 936
rect 578 813 581 943
rect 586 943 605 946
rect 586 913 589 943
rect 586 823 589 906
rect 602 903 605 926
rect 594 786 597 816
rect 610 793 613 806
rect 586 783 597 786
rect 586 726 589 783
rect 602 733 605 786
rect 538 703 541 726
rect 546 716 549 726
rect 586 723 597 726
rect 546 713 557 716
rect 514 693 525 696
rect 498 683 509 686
rect 490 613 493 636
rect 498 606 501 683
rect 506 613 509 646
rect 522 636 525 693
rect 514 633 525 636
rect 514 613 517 633
rect 498 603 525 606
rect 458 543 469 546
rect 458 523 461 543
rect 482 533 485 546
rect 498 523 501 596
rect 434 443 453 446
rect 362 403 365 416
rect 370 413 381 416
rect 338 356 341 376
rect 338 353 349 356
rect 290 316 293 323
rect 322 316 325 346
rect 282 313 293 316
rect 306 313 325 316
rect 282 213 285 313
rect 330 303 333 326
rect 346 266 349 353
rect 370 333 373 413
rect 378 383 381 406
rect 410 316 413 336
rect 330 263 349 266
rect 402 313 413 316
rect 402 266 405 313
rect 402 263 413 266
rect 306 193 309 206
rect 330 193 333 263
rect 378 193 381 216
rect 410 213 413 263
rect 418 206 421 326
rect 426 303 429 336
rect 434 323 437 443
rect 442 336 445 416
rect 466 403 469 416
rect 482 413 485 516
rect 506 496 509 586
rect 522 533 525 603
rect 554 566 557 713
rect 594 703 597 723
rect 618 713 621 916
rect 626 913 629 926
rect 634 846 637 1003
rect 642 996 645 1016
rect 650 1003 653 1016
rect 642 993 649 996
rect 646 936 649 993
rect 658 943 661 1006
rect 666 986 669 1076
rect 674 1013 677 1026
rect 666 983 673 986
rect 670 936 673 983
rect 646 933 653 936
rect 626 843 637 846
rect 610 623 613 706
rect 570 593 573 616
rect 594 603 597 616
rect 610 593 613 606
rect 554 563 573 566
rect 490 493 509 496
rect 442 333 461 336
rect 490 333 493 493
rect 514 473 517 526
rect 498 313 501 416
rect 506 383 509 406
rect 514 393 517 416
rect 522 413 525 516
rect 530 493 533 526
rect 522 323 525 406
rect 530 333 533 406
rect 538 343 541 416
rect 546 413 549 546
rect 570 426 573 563
rect 578 513 581 586
rect 626 583 629 843
rect 634 723 637 816
rect 642 803 645 826
rect 642 733 645 796
rect 650 773 653 933
rect 666 933 673 936
rect 682 933 685 1153
rect 730 1123 733 1136
rect 738 1133 741 1153
rect 738 1113 741 1126
rect 666 843 669 933
rect 666 813 669 836
rect 674 793 677 896
rect 682 813 685 916
rect 690 886 693 1016
rect 698 966 701 1026
rect 706 983 709 1006
rect 698 963 709 966
rect 698 933 701 956
rect 698 896 701 926
rect 706 923 709 963
rect 714 953 717 1046
rect 722 956 725 1006
rect 730 1003 733 1096
rect 746 1073 749 1146
rect 754 1133 757 1153
rect 762 1133 765 1146
rect 754 1123 765 1126
rect 754 1013 757 1066
rect 786 1056 789 1126
rect 810 1093 813 1576
rect 826 1563 829 1656
rect 834 1583 837 1616
rect 850 1613 853 1783
rect 858 1733 861 1793
rect 906 1756 909 1936
rect 922 1933 925 1993
rect 954 1923 957 1956
rect 914 1803 917 1816
rect 906 1753 913 1756
rect 858 1713 861 1726
rect 910 1706 913 1753
rect 906 1703 913 1706
rect 906 1653 909 1703
rect 922 1653 925 1786
rect 842 1593 845 1606
rect 818 1533 821 1556
rect 850 1553 853 1606
rect 858 1596 861 1616
rect 866 1603 869 1616
rect 874 1596 877 1606
rect 858 1593 877 1596
rect 882 1593 885 1616
rect 890 1613 893 1626
rect 906 1603 909 1636
rect 930 1633 933 1866
rect 938 1723 941 1736
rect 930 1613 933 1626
rect 826 1543 845 1546
rect 818 1363 821 1526
rect 826 1523 829 1543
rect 834 1526 837 1536
rect 842 1533 845 1543
rect 834 1523 845 1526
rect 826 1286 829 1426
rect 818 1283 829 1286
rect 818 1133 821 1283
rect 834 1253 837 1516
rect 842 1433 845 1523
rect 850 1503 853 1526
rect 858 1513 861 1526
rect 842 1323 845 1416
rect 850 1413 853 1486
rect 850 1393 853 1406
rect 858 1346 861 1436
rect 866 1363 869 1456
rect 850 1343 861 1346
rect 850 1246 853 1343
rect 842 1243 853 1246
rect 842 1203 845 1236
rect 874 1233 877 1536
rect 898 1533 901 1556
rect 898 1513 901 1526
rect 906 1496 909 1596
rect 894 1493 909 1496
rect 882 1363 885 1446
rect 894 1436 897 1493
rect 914 1453 917 1516
rect 890 1433 897 1436
rect 922 1433 925 1566
rect 938 1513 941 1656
rect 946 1496 949 1776
rect 962 1773 965 1946
rect 970 1903 973 2116
rect 994 2043 997 2156
rect 994 2016 997 2026
rect 978 2013 989 2016
rect 994 2013 1005 2016
rect 978 1933 981 2013
rect 994 1993 997 2006
rect 1002 1986 1005 2013
rect 994 1983 1005 1986
rect 994 1923 997 1983
rect 1010 1963 1013 2056
rect 1018 2003 1021 2206
rect 1026 2196 1029 2213
rect 1026 2193 1033 2196
rect 1042 2193 1045 2206
rect 1030 2046 1033 2193
rect 1058 2153 1061 2253
rect 1082 2193 1085 2216
rect 1042 2123 1045 2136
rect 1074 2133 1085 2136
rect 1026 2043 1033 2046
rect 1026 2013 1029 2043
rect 1042 2013 1045 2116
rect 1074 2106 1077 2126
rect 1098 2123 1101 2393
rect 1138 2213 1141 2336
rect 1146 2213 1149 2476
rect 1162 2413 1165 2426
rect 1162 2333 1165 2406
rect 1170 2326 1173 2526
rect 1178 2523 1197 2526
rect 1186 2506 1189 2523
rect 1182 2503 1189 2506
rect 1182 2436 1185 2503
rect 1194 2443 1197 2516
rect 1202 2436 1205 2496
rect 1182 2433 1189 2436
rect 1186 2416 1189 2433
rect 1194 2433 1205 2436
rect 1194 2423 1197 2433
rect 1186 2413 1197 2416
rect 1202 2413 1205 2433
rect 1178 2403 1189 2406
rect 1162 2323 1173 2326
rect 1162 2246 1165 2323
rect 1154 2243 1165 2246
rect 1154 2213 1157 2243
rect 1170 2223 1189 2226
rect 1138 2203 1149 2206
rect 1146 2173 1149 2203
rect 1170 2193 1173 2206
rect 1178 2136 1181 2216
rect 1106 2123 1109 2136
rect 1066 2103 1077 2106
rect 1066 2046 1069 2103
rect 1066 2043 1077 2046
rect 1026 1943 1029 2006
rect 1074 2003 1077 2043
rect 1082 2013 1085 2116
rect 1034 1946 1037 1966
rect 1090 1956 1093 2066
rect 1114 2053 1117 2136
rect 1162 2133 1181 2136
rect 1138 2083 1141 2126
rect 1098 2023 1101 2036
rect 1082 1953 1093 1956
rect 1034 1943 1045 1946
rect 994 1903 997 1916
rect 1010 1863 1013 1936
rect 1042 1896 1045 1943
rect 1082 1936 1085 1953
rect 1078 1933 1085 1936
rect 1034 1893 1045 1896
rect 978 1813 981 1826
rect 994 1733 997 1806
rect 1010 1803 1013 1816
rect 1018 1813 1021 1826
rect 1034 1786 1037 1893
rect 1058 1813 1061 1926
rect 1078 1886 1081 1933
rect 1090 1896 1093 1946
rect 1098 1933 1101 2006
rect 1106 1963 1109 2026
rect 1154 2003 1157 2016
rect 1162 2003 1165 2133
rect 1186 2123 1189 2223
rect 1194 2123 1197 2413
rect 1210 2403 1213 2426
rect 1210 2203 1213 2216
rect 1202 2123 1205 2136
rect 1186 2043 1189 2116
rect 1210 2083 1213 2196
rect 1218 2063 1221 2406
rect 1226 2376 1229 2536
rect 1250 2523 1253 2546
rect 1250 2413 1253 2456
rect 1274 2413 1277 2446
rect 1282 2403 1285 2426
rect 1290 2413 1293 2426
rect 1306 2403 1309 2546
rect 1322 2533 1325 2556
rect 1330 2533 1333 2586
rect 1346 2553 1349 2637
rect 1314 2396 1317 2416
rect 1322 2413 1325 2426
rect 1306 2393 1317 2396
rect 1226 2373 1245 2376
rect 1242 2266 1245 2373
rect 1226 2263 1245 2266
rect 1178 2013 1181 2036
rect 1186 2013 1189 2026
rect 1210 1983 1213 2006
rect 1226 2003 1229 2263
rect 1234 2116 1237 2216
rect 1258 2203 1261 2226
rect 1282 2213 1285 2376
rect 1306 2313 1309 2393
rect 1330 2373 1333 2526
rect 1354 2503 1357 2526
rect 1378 2513 1381 2556
rect 1386 2483 1389 2536
rect 1434 2533 1437 2546
rect 1442 2533 1445 2556
rect 1490 2533 1493 2546
rect 1410 2513 1413 2526
rect 1370 2413 1373 2436
rect 1338 2383 1341 2406
rect 1346 2363 1349 2406
rect 1314 2333 1317 2346
rect 1330 2286 1333 2336
rect 1354 2323 1357 2346
rect 1394 2333 1397 2406
rect 1418 2403 1421 2426
rect 1410 2323 1413 2386
rect 1426 2373 1429 2416
rect 1450 2413 1453 2446
rect 1466 2436 1469 2526
rect 1530 2466 1533 2526
rect 1530 2463 1541 2466
rect 1466 2433 1485 2436
rect 1474 2376 1477 2406
rect 1466 2373 1477 2376
rect 1418 2323 1421 2336
rect 1330 2283 1341 2286
rect 1418 2283 1421 2316
rect 1442 2313 1445 2326
rect 1466 2303 1469 2373
rect 1306 2213 1309 2226
rect 1274 2173 1277 2206
rect 1306 2203 1317 2206
rect 1322 2186 1325 2206
rect 1338 2203 1341 2283
rect 1474 2226 1477 2346
rect 1482 2233 1485 2433
rect 1490 2343 1493 2416
rect 1538 2403 1541 2463
rect 1546 2413 1549 2536
rect 1554 2473 1557 2536
rect 1578 2493 1581 2526
rect 1602 2523 1605 2536
rect 1634 2513 1637 2526
rect 1570 2413 1573 2426
rect 1498 2256 1501 2376
rect 1546 2356 1549 2406
rect 1594 2383 1597 2406
rect 1602 2403 1605 2446
rect 1658 2436 1661 2536
rect 1714 2533 1717 2546
rect 1802 2543 1829 2546
rect 1690 2483 1693 2526
rect 1698 2493 1701 2526
rect 1722 2523 1725 2536
rect 1658 2433 1669 2436
rect 1618 2373 1621 2426
rect 1642 2413 1645 2426
rect 1666 2403 1669 2433
rect 1674 2403 1677 2426
rect 1706 2413 1709 2426
rect 1546 2353 1565 2356
rect 1554 2333 1557 2346
rect 1562 2333 1565 2353
rect 1570 2343 1581 2346
rect 1490 2253 1501 2256
rect 1362 2203 1365 2216
rect 1322 2183 1333 2186
rect 1242 2126 1245 2136
rect 1242 2123 1253 2126
rect 1234 2113 1245 2116
rect 1242 2093 1245 2113
rect 1250 2013 1253 2123
rect 1266 2076 1269 2106
rect 1274 2093 1277 2136
rect 1282 2133 1285 2156
rect 1330 2133 1333 2183
rect 1266 2073 1273 2076
rect 1146 1933 1149 1966
rect 1146 1913 1149 1926
rect 1162 1903 1165 1936
rect 1090 1893 1101 1896
rect 1078 1883 1085 1886
rect 1018 1783 1037 1786
rect 954 1563 957 1666
rect 970 1553 973 1726
rect 978 1713 981 1726
rect 978 1613 989 1616
rect 978 1593 981 1613
rect 986 1603 997 1606
rect 1002 1576 1005 1736
rect 986 1573 1005 1576
rect 962 1533 965 1546
rect 970 1533 981 1536
rect 954 1503 957 1526
rect 938 1493 949 1496
rect 938 1443 941 1493
rect 890 1373 893 1433
rect 914 1423 933 1426
rect 898 1396 901 1416
rect 906 1403 909 1416
rect 914 1413 917 1423
rect 914 1396 917 1406
rect 898 1393 917 1396
rect 898 1333 901 1346
rect 922 1323 925 1416
rect 930 1393 933 1423
rect 946 1343 949 1486
rect 970 1413 973 1526
rect 978 1493 981 1526
rect 978 1406 981 1436
rect 970 1403 981 1406
rect 970 1396 973 1403
rect 966 1393 973 1396
rect 966 1286 969 1393
rect 962 1283 969 1286
rect 882 1213 885 1226
rect 850 1153 853 1186
rect 858 1163 861 1206
rect 882 1156 885 1186
rect 906 1173 909 1226
rect 914 1213 917 1236
rect 938 1213 941 1226
rect 946 1213 949 1256
rect 962 1213 965 1283
rect 978 1253 981 1396
rect 986 1353 989 1573
rect 994 1523 997 1546
rect 1002 1523 1005 1536
rect 1010 1533 1013 1616
rect 1018 1573 1021 1783
rect 1034 1733 1037 1756
rect 1042 1723 1045 1806
rect 1042 1696 1045 1716
rect 1034 1693 1045 1696
rect 1034 1646 1037 1693
rect 1034 1643 1045 1646
rect 1026 1613 1029 1626
rect 994 1343 997 1416
rect 994 1313 997 1336
rect 874 1153 885 1156
rect 874 1136 877 1153
rect 866 1133 877 1136
rect 882 1133 885 1146
rect 786 1053 805 1056
rect 778 1003 781 1036
rect 786 1013 789 1046
rect 802 1013 805 1053
rect 818 1013 821 1126
rect 722 953 733 956
rect 722 933 725 946
rect 722 913 725 926
rect 698 893 717 896
rect 690 883 709 886
rect 690 823 693 836
rect 682 783 685 806
rect 698 776 701 826
rect 706 813 709 883
rect 714 803 717 893
rect 722 813 725 826
rect 730 806 733 953
rect 738 813 741 846
rect 722 803 733 806
rect 642 706 645 726
rect 674 716 677 736
rect 666 713 677 716
rect 642 703 653 706
rect 650 646 653 703
rect 642 643 653 646
rect 666 646 669 713
rect 666 643 677 646
rect 634 603 637 626
rect 642 613 645 643
rect 666 616 669 626
rect 650 596 653 616
rect 642 593 653 596
rect 658 613 669 616
rect 674 613 677 643
rect 562 423 573 426
rect 546 366 549 406
rect 554 373 557 416
rect 578 413 581 436
rect 562 383 565 406
rect 546 363 557 366
rect 570 363 573 406
rect 586 366 589 566
rect 594 523 597 546
rect 610 523 629 526
rect 610 506 613 523
rect 610 503 621 506
rect 578 363 589 366
rect 594 363 597 406
rect 602 376 605 486
rect 618 446 621 503
rect 634 483 637 536
rect 642 523 645 593
rect 658 583 661 613
rect 666 603 677 606
rect 658 533 661 546
rect 666 526 669 536
rect 666 523 677 526
rect 666 503 669 516
rect 674 483 677 523
rect 682 476 685 776
rect 690 773 701 776
rect 690 733 693 773
rect 746 733 749 976
rect 762 933 765 986
rect 770 943 773 956
rect 778 936 781 996
rect 786 943 789 1006
rect 834 1003 837 1116
rect 842 1103 845 1126
rect 866 1113 869 1133
rect 842 1003 845 1096
rect 866 1013 869 1026
rect 874 1013 877 1126
rect 890 1113 893 1166
rect 954 1156 957 1176
rect 950 1153 957 1156
rect 914 1113 917 1126
rect 938 1123 941 1146
rect 950 1066 953 1153
rect 962 1133 965 1206
rect 970 1133 973 1156
rect 950 1063 957 1066
rect 890 1003 893 1016
rect 898 1003 901 1036
rect 946 1013 949 1046
rect 802 956 805 986
rect 794 953 805 956
rect 778 933 789 936
rect 778 893 781 916
rect 754 786 757 816
rect 762 803 765 856
rect 786 833 789 933
rect 794 823 797 953
rect 802 903 805 946
rect 810 933 813 956
rect 810 843 813 916
rect 754 783 761 786
rect 758 726 761 783
rect 706 603 709 616
rect 714 596 717 726
rect 754 723 761 726
rect 754 613 757 723
rect 770 613 773 786
rect 690 533 693 596
rect 706 593 717 596
rect 706 576 709 593
rect 698 573 709 576
rect 738 576 741 596
rect 754 586 757 606
rect 754 583 765 586
rect 738 573 757 576
rect 690 516 693 526
rect 698 523 701 573
rect 706 523 717 526
rect 690 513 717 516
rect 722 513 725 566
rect 610 443 621 446
rect 666 473 685 476
rect 610 403 613 443
rect 602 373 613 376
rect 554 356 557 363
rect 578 356 581 363
rect 554 353 581 356
rect 554 333 557 353
rect 426 213 429 296
rect 442 223 445 266
rect 546 263 549 326
rect 562 263 565 326
rect 562 216 565 226
rect 402 203 421 206
rect 250 173 269 176
rect 226 133 229 146
rect 202 -147 205 126
rect 210 123 229 126
rect 250 123 253 173
rect 258 133 261 166
rect 274 133 277 156
rect 322 123 325 146
rect 378 133 381 146
rect 226 113 229 123
rect 290 -141 293 96
rect 354 93 357 126
rect 378 113 381 126
rect 402 123 405 203
rect 442 193 445 206
rect 410 133 413 166
rect 426 133 429 156
rect 450 136 453 216
rect 506 193 509 216
rect 554 213 565 216
rect 530 153 533 206
rect 546 183 549 206
rect 450 133 461 136
rect 458 76 461 133
rect 474 123 477 146
rect 530 133 533 146
rect 450 73 461 76
rect 450 16 453 73
rect 450 13 461 16
rect 458 -135 461 13
rect 474 -125 477 116
rect 506 113 509 126
rect 530 113 533 126
rect 554 123 557 213
rect 562 193 565 206
rect 562 133 565 166
rect 578 133 581 346
rect 610 296 613 373
rect 626 353 629 406
rect 666 383 669 473
rect 674 403 677 416
rect 626 323 629 346
rect 682 333 685 346
rect 690 326 693 506
rect 698 416 701 486
rect 714 423 717 513
rect 730 496 733 526
rect 726 493 733 496
rect 698 413 709 416
rect 698 386 701 413
rect 706 403 717 406
rect 698 383 705 386
rect 594 293 613 296
rect 594 213 597 293
rect 594 143 597 206
rect 610 163 613 206
rect 642 166 645 286
rect 666 256 669 326
rect 682 323 693 326
rect 682 276 685 323
rect 702 306 705 383
rect 726 346 729 493
rect 738 413 741 526
rect 746 516 749 536
rect 754 533 757 573
rect 762 553 765 583
rect 762 533 765 546
rect 770 523 773 576
rect 778 563 781 656
rect 746 513 757 516
rect 778 513 781 536
rect 786 533 789 606
rect 794 603 797 776
rect 810 693 813 836
rect 818 813 821 826
rect 826 773 829 966
rect 842 933 845 996
rect 842 896 845 926
rect 842 893 853 896
rect 850 826 853 893
rect 890 833 893 936
rect 898 933 901 986
rect 946 943 949 1006
rect 954 963 957 1063
rect 846 823 853 826
rect 834 736 837 816
rect 846 756 849 823
rect 826 733 837 736
rect 842 753 849 756
rect 826 713 829 733
rect 842 703 845 753
rect 818 613 821 626
rect 850 613 853 736
rect 858 716 861 806
rect 866 723 869 806
rect 898 803 901 816
rect 882 723 885 746
rect 858 713 877 716
rect 842 593 845 606
rect 802 583 813 586
rect 794 533 797 576
rect 802 533 805 546
rect 754 436 757 513
rect 786 436 789 526
rect 746 433 757 436
rect 782 433 789 436
rect 746 413 749 433
rect 726 343 733 346
rect 714 323 717 336
rect 730 323 733 343
rect 698 303 705 306
rect 698 283 701 303
rect 682 273 701 276
rect 666 253 677 256
rect 674 226 677 253
rect 674 223 685 226
rect 658 193 661 216
rect 642 163 649 166
rect 562 113 565 126
rect 626 123 629 146
rect 646 96 649 163
rect 642 93 649 96
rect 642 76 645 93
rect 634 73 645 76
rect 634 16 637 73
rect 634 13 645 16
rect 642 -116 645 13
rect 658 -106 661 186
rect 682 176 685 223
rect 690 183 693 216
rect 682 173 693 176
rect 682 133 685 146
rect 666 96 669 126
rect 682 113 685 126
rect 690 106 693 173
rect 698 123 701 273
rect 738 206 741 406
rect 782 376 785 433
rect 802 426 805 526
rect 810 523 813 583
rect 818 513 821 536
rect 826 533 829 546
rect 794 423 805 426
rect 794 376 797 423
rect 802 383 805 416
rect 826 413 829 526
rect 834 523 837 586
rect 850 573 853 606
rect 858 583 861 706
rect 874 613 877 626
rect 890 613 893 636
rect 898 613 901 756
rect 906 713 909 826
rect 914 753 917 926
rect 922 813 925 826
rect 866 593 869 606
rect 874 586 877 606
rect 882 593 885 606
rect 866 583 877 586
rect 898 586 901 606
rect 906 603 909 626
rect 914 596 917 726
rect 906 593 917 596
rect 922 586 925 726
rect 930 716 933 836
rect 938 823 941 836
rect 946 723 949 926
rect 954 823 957 936
rect 962 923 965 1126
rect 978 1116 981 1246
rect 1002 1213 1005 1326
rect 1010 1203 1013 1476
rect 1018 1323 1021 1556
rect 1026 1523 1029 1606
rect 1026 1366 1029 1516
rect 1034 1413 1037 1616
rect 1042 1603 1045 1643
rect 1050 1613 1053 1736
rect 1042 1493 1045 1576
rect 1058 1553 1061 1806
rect 1082 1783 1085 1883
rect 1098 1826 1101 1893
rect 1186 1876 1189 1956
rect 1234 1946 1237 1966
rect 1258 1953 1261 2056
rect 1270 1986 1273 2073
rect 1298 2043 1301 2126
rect 1266 1983 1273 1986
rect 1266 1963 1269 1983
rect 1230 1943 1237 1946
rect 1090 1823 1101 1826
rect 1178 1873 1189 1876
rect 1066 1723 1069 1746
rect 1074 1733 1077 1756
rect 1090 1716 1093 1823
rect 1178 1806 1181 1873
rect 1202 1813 1205 1926
rect 1210 1876 1213 1906
rect 1230 1886 1233 1943
rect 1242 1896 1245 1926
rect 1250 1923 1253 1936
rect 1298 1933 1301 2036
rect 1306 2013 1309 2096
rect 1338 2053 1341 2136
rect 1362 2073 1365 2126
rect 1386 2066 1389 2156
rect 1418 2153 1421 2216
rect 1394 2103 1397 2136
rect 1418 2083 1421 2126
rect 1442 2106 1445 2136
rect 1426 2103 1445 2106
rect 1370 2063 1389 2066
rect 1338 2013 1341 2036
rect 1306 2003 1317 2006
rect 1362 2003 1365 2026
rect 1370 2003 1373 2063
rect 1394 2013 1397 2036
rect 1418 2013 1421 2066
rect 1418 1986 1421 2006
rect 1426 2003 1429 2103
rect 1442 2023 1445 2056
rect 1450 2043 1453 2126
rect 1458 2116 1461 2226
rect 1474 2223 1485 2226
rect 1482 2143 1485 2223
rect 1490 2186 1493 2253
rect 1498 2193 1501 2236
rect 1490 2183 1501 2186
rect 1498 2123 1501 2183
rect 1506 2133 1509 2156
rect 1458 2113 1469 2116
rect 1466 2093 1469 2106
rect 1482 2103 1485 2116
rect 1458 2013 1461 2026
rect 1306 1933 1309 1986
rect 1354 1933 1357 1986
rect 1410 1983 1421 1986
rect 1362 1933 1365 1956
rect 1306 1913 1309 1926
rect 1242 1893 1261 1896
rect 1230 1883 1237 1886
rect 1210 1873 1221 1876
rect 1218 1806 1221 1873
rect 1098 1723 1101 1806
rect 1106 1723 1109 1736
rect 1114 1733 1117 1756
rect 1114 1716 1117 1726
rect 1122 1723 1125 1736
rect 1090 1713 1117 1716
rect 1106 1613 1109 1636
rect 1050 1513 1053 1526
rect 1066 1483 1069 1536
rect 1090 1513 1093 1526
rect 1050 1413 1053 1426
rect 1034 1383 1037 1406
rect 1082 1403 1085 1456
rect 1026 1363 1037 1366
rect 1026 1333 1029 1356
rect 1034 1333 1037 1363
rect 1034 1313 1037 1326
rect 1010 1163 1013 1196
rect 1018 1173 1021 1266
rect 974 1113 981 1116
rect 974 1026 977 1113
rect 970 1023 977 1026
rect 970 1003 973 1023
rect 1002 1013 1005 1026
rect 978 913 981 1006
rect 1026 1003 1029 1256
rect 1034 1153 1037 1166
rect 994 923 1005 926
rect 994 903 997 916
rect 1002 903 1005 916
rect 1010 913 1013 946
rect 1018 923 1029 926
rect 1034 853 1037 1146
rect 1042 993 1045 1366
rect 1066 1333 1069 1346
rect 1074 1333 1077 1356
rect 1050 1143 1053 1256
rect 1058 1163 1061 1326
rect 1082 1323 1085 1396
rect 1066 1213 1069 1276
rect 1082 1223 1085 1296
rect 1090 1253 1093 1496
rect 1098 1436 1101 1576
rect 1106 1443 1109 1606
rect 1114 1523 1117 1713
rect 1122 1563 1125 1626
rect 1130 1586 1133 1726
rect 1138 1706 1141 1736
rect 1146 1723 1149 1806
rect 1178 1803 1189 1806
rect 1154 1723 1157 1736
rect 1138 1703 1149 1706
rect 1162 1703 1165 1726
rect 1146 1636 1149 1703
rect 1170 1696 1173 1736
rect 1138 1633 1149 1636
rect 1162 1693 1173 1696
rect 1138 1603 1141 1633
rect 1146 1596 1149 1616
rect 1162 1613 1165 1693
rect 1170 1603 1173 1616
rect 1146 1593 1157 1596
rect 1130 1583 1137 1586
rect 1134 1506 1137 1583
rect 1130 1503 1137 1506
rect 1130 1486 1133 1503
rect 1122 1483 1133 1486
rect 1146 1483 1149 1566
rect 1154 1533 1157 1593
rect 1178 1563 1181 1706
rect 1186 1623 1189 1803
rect 1210 1803 1221 1806
rect 1210 1733 1213 1803
rect 1234 1733 1237 1883
rect 1258 1776 1261 1893
rect 1242 1773 1261 1776
rect 1194 1713 1197 1726
rect 1210 1706 1213 1726
rect 1234 1713 1237 1726
rect 1194 1703 1213 1706
rect 1242 1703 1245 1773
rect 1186 1583 1189 1616
rect 1194 1596 1197 1703
rect 1202 1603 1205 1636
rect 1290 1633 1293 1766
rect 1298 1733 1301 1746
rect 1250 1596 1253 1606
rect 1258 1603 1261 1616
rect 1266 1613 1269 1626
rect 1266 1603 1277 1606
rect 1266 1596 1269 1603
rect 1194 1593 1205 1596
rect 1250 1593 1269 1596
rect 1202 1533 1205 1593
rect 1210 1533 1213 1566
rect 1098 1433 1109 1436
rect 1106 1423 1109 1433
rect 1122 1413 1125 1483
rect 1138 1413 1141 1426
rect 1146 1413 1149 1436
rect 1162 1423 1165 1506
rect 1170 1413 1173 1526
rect 1178 1466 1181 1526
rect 1202 1473 1205 1526
rect 1178 1463 1197 1466
rect 1194 1413 1197 1463
rect 1138 1393 1141 1406
rect 1146 1386 1149 1406
rect 1202 1403 1205 1416
rect 1218 1413 1237 1416
rect 1146 1383 1173 1386
rect 1098 1356 1101 1376
rect 1098 1353 1105 1356
rect 1102 1246 1105 1353
rect 1122 1333 1125 1346
rect 1130 1333 1133 1356
rect 1114 1256 1117 1326
rect 1146 1273 1149 1326
rect 1154 1323 1157 1376
rect 1162 1373 1173 1376
rect 1162 1263 1165 1373
rect 1170 1326 1173 1366
rect 1178 1333 1181 1356
rect 1194 1333 1197 1346
rect 1170 1323 1177 1326
rect 1114 1253 1125 1256
rect 1098 1243 1105 1246
rect 1090 1213 1093 1236
rect 1098 1213 1101 1243
rect 1122 1213 1125 1253
rect 1174 1246 1177 1323
rect 1186 1263 1189 1326
rect 1202 1306 1205 1396
rect 1210 1353 1213 1406
rect 1226 1356 1229 1406
rect 1234 1403 1237 1413
rect 1242 1363 1245 1446
rect 1258 1426 1261 1546
rect 1266 1513 1269 1526
rect 1250 1423 1261 1426
rect 1274 1423 1277 1566
rect 1282 1543 1285 1616
rect 1290 1556 1293 1616
rect 1298 1613 1301 1626
rect 1298 1593 1301 1606
rect 1306 1563 1309 1876
rect 1330 1826 1333 1926
rect 1338 1913 1341 1926
rect 1386 1906 1389 1926
rect 1378 1903 1389 1906
rect 1378 1856 1381 1903
rect 1378 1853 1389 1856
rect 1322 1823 1333 1826
rect 1370 1823 1373 1836
rect 1386 1826 1389 1853
rect 1394 1846 1397 1946
rect 1394 1843 1405 1846
rect 1378 1823 1389 1826
rect 1322 1766 1325 1823
rect 1322 1763 1333 1766
rect 1314 1743 1325 1746
rect 1314 1723 1317 1736
rect 1322 1723 1325 1743
rect 1330 1733 1333 1763
rect 1330 1703 1333 1726
rect 1338 1723 1341 1816
rect 1354 1643 1357 1726
rect 1362 1723 1365 1736
rect 1378 1733 1381 1823
rect 1402 1786 1405 1843
rect 1410 1836 1413 1983
rect 1474 1946 1477 2036
rect 1482 2016 1485 2096
rect 1490 2053 1493 2116
rect 1514 2113 1517 2126
rect 1522 2076 1525 2216
rect 1530 2173 1533 2326
rect 1570 2286 1573 2343
rect 1562 2283 1573 2286
rect 1538 2133 1541 2236
rect 1546 2196 1549 2216
rect 1562 2213 1565 2283
rect 1578 2206 1581 2336
rect 1586 2273 1589 2336
rect 1586 2213 1589 2236
rect 1546 2193 1557 2196
rect 1554 2133 1557 2193
rect 1562 2153 1565 2206
rect 1570 2193 1573 2206
rect 1578 2203 1589 2206
rect 1594 2203 1597 2306
rect 1610 2293 1613 2326
rect 1634 2303 1637 2386
rect 1642 2333 1645 2376
rect 1698 2343 1701 2356
rect 1722 2336 1725 2516
rect 1770 2493 1773 2526
rect 1778 2513 1781 2536
rect 1802 2533 1805 2543
rect 1810 2533 1829 2536
rect 1850 2533 1853 2546
rect 1866 2533 1893 2536
rect 1906 2533 1909 2546
rect 2002 2543 2021 2546
rect 1762 2433 1765 2456
rect 1730 2353 1733 2406
rect 1754 2396 1757 2426
rect 1738 2393 1757 2396
rect 1778 2406 1781 2466
rect 1786 2423 1789 2526
rect 1794 2413 1797 2496
rect 1810 2443 1813 2526
rect 1818 2453 1821 2533
rect 1842 2493 1845 2526
rect 1858 2463 1861 2516
rect 1866 2513 1869 2533
rect 1882 2513 1885 2526
rect 1890 2506 1893 2526
rect 1890 2503 1901 2506
rect 1810 2423 1813 2436
rect 1818 2413 1821 2426
rect 1842 2423 1845 2436
rect 1850 2413 1853 2446
rect 1778 2403 1821 2406
rect 1586 2146 1589 2203
rect 1642 2193 1645 2206
rect 1562 2143 1573 2146
rect 1586 2143 1605 2146
rect 1530 2113 1533 2126
rect 1538 2093 1541 2126
rect 1522 2073 1533 2076
rect 1490 2023 1493 2036
rect 1498 2023 1501 2036
rect 1482 2013 1493 2016
rect 1506 1996 1509 2026
rect 1514 2023 1517 2036
rect 1522 2006 1525 2056
rect 1530 2013 1533 2073
rect 1538 2033 1549 2036
rect 1470 1943 1477 1946
rect 1498 1993 1509 1996
rect 1410 1833 1421 1836
rect 1410 1796 1413 1826
rect 1418 1803 1421 1833
rect 1410 1793 1421 1796
rect 1402 1783 1413 1786
rect 1378 1723 1389 1726
rect 1290 1553 1301 1556
rect 1290 1423 1293 1536
rect 1298 1523 1301 1553
rect 1306 1533 1309 1546
rect 1314 1493 1317 1626
rect 1338 1613 1341 1626
rect 1394 1616 1397 1736
rect 1410 1713 1413 1783
rect 1418 1733 1421 1793
rect 1426 1783 1429 1816
rect 1434 1813 1437 1926
rect 1434 1793 1437 1806
rect 1442 1803 1445 1826
rect 1442 1716 1445 1736
rect 1450 1723 1453 1816
rect 1458 1803 1461 1926
rect 1470 1846 1473 1943
rect 1470 1843 1477 1846
rect 1442 1713 1453 1716
rect 1458 1713 1461 1726
rect 1466 1723 1469 1816
rect 1474 1813 1477 1843
rect 1482 1803 1485 1936
rect 1498 1873 1501 1993
rect 1506 1866 1509 1916
rect 1514 1896 1517 2006
rect 1522 2003 1533 2006
rect 1538 2003 1541 2026
rect 1530 1913 1533 2003
rect 1546 1926 1549 2033
rect 1554 2013 1557 2116
rect 1562 2053 1565 2143
rect 1570 2113 1573 2126
rect 1562 2013 1565 2046
rect 1586 2033 1589 2126
rect 1578 2013 1581 2026
rect 1570 1983 1573 2006
rect 1586 1976 1589 2006
rect 1578 1973 1589 1976
rect 1538 1923 1549 1926
rect 1554 1923 1557 1936
rect 1562 1913 1565 1926
rect 1514 1893 1525 1896
rect 1498 1863 1509 1866
rect 1490 1813 1493 1826
rect 1482 1723 1485 1786
rect 1498 1783 1501 1863
rect 1506 1793 1509 1816
rect 1514 1803 1517 1816
rect 1506 1726 1509 1736
rect 1490 1723 1509 1726
rect 1514 1723 1517 1796
rect 1522 1773 1525 1893
rect 1570 1846 1573 1936
rect 1578 1923 1581 1973
rect 1594 1966 1597 2126
rect 1602 2123 1605 2143
rect 1610 2056 1613 2166
rect 1586 1963 1597 1966
rect 1602 2053 1613 2056
rect 1586 1933 1589 1963
rect 1602 1933 1605 2053
rect 1610 1986 1613 2036
rect 1618 1993 1621 2006
rect 1610 1983 1621 1986
rect 1626 1983 1629 2156
rect 1650 2153 1653 2216
rect 1634 2113 1637 2136
rect 1642 2123 1645 2146
rect 1650 2033 1653 2136
rect 1658 2123 1661 2326
rect 1666 2303 1669 2336
rect 1722 2333 1733 2336
rect 1738 2326 1741 2393
rect 1682 2236 1685 2326
rect 1722 2323 1741 2326
rect 1722 2306 1725 2323
rect 1714 2303 1725 2306
rect 1714 2246 1717 2303
rect 1714 2243 1725 2246
rect 1678 2233 1685 2236
rect 1666 2163 1669 2206
rect 1678 2166 1681 2233
rect 1722 2226 1725 2243
rect 1678 2163 1685 2166
rect 1666 2133 1669 2156
rect 1674 2133 1677 2146
rect 1666 2113 1669 2126
rect 1682 2123 1685 2163
rect 1690 2133 1693 2226
rect 1714 2223 1725 2226
rect 1730 2216 1733 2316
rect 1698 2133 1701 2206
rect 1714 2203 1717 2216
rect 1722 2213 1733 2216
rect 1714 2133 1717 2176
rect 1738 2146 1741 2196
rect 1746 2193 1749 2336
rect 1762 2323 1765 2356
rect 1738 2143 1749 2146
rect 1706 2103 1709 2126
rect 1746 2123 1749 2143
rect 1754 2133 1757 2316
rect 1762 2193 1765 2216
rect 1770 2213 1773 2336
rect 1778 2293 1781 2403
rect 1858 2373 1861 2406
rect 1794 2353 1813 2356
rect 1786 2226 1789 2326
rect 1794 2296 1797 2353
rect 1802 2333 1805 2346
rect 1810 2333 1813 2353
rect 1818 2336 1821 2346
rect 1834 2343 1837 2366
rect 1866 2343 1869 2426
rect 1874 2403 1877 2496
rect 1898 2426 1901 2503
rect 1890 2423 1901 2426
rect 1818 2333 1829 2336
rect 1810 2306 1813 2326
rect 1818 2323 1821 2333
rect 1810 2303 1817 2306
rect 1794 2293 1805 2296
rect 1778 2223 1789 2226
rect 1770 2186 1773 2206
rect 1762 2183 1773 2186
rect 1762 2133 1765 2183
rect 1778 2123 1781 2223
rect 1786 2203 1789 2216
rect 1762 2096 1765 2116
rect 1754 2093 1765 2096
rect 1706 2016 1709 2036
rect 1618 1926 1621 1983
rect 1634 1933 1637 2016
rect 1642 2003 1645 2016
rect 1706 2013 1713 2016
rect 1642 1926 1645 1966
rect 1690 1933 1693 2006
rect 1594 1913 1597 1926
rect 1570 1843 1581 1846
rect 1562 1823 1565 1836
rect 1570 1823 1573 1836
rect 1538 1813 1573 1816
rect 1466 1713 1477 1716
rect 1466 1703 1469 1713
rect 1482 1703 1485 1716
rect 1490 1703 1493 1723
rect 1322 1533 1333 1536
rect 1338 1533 1341 1546
rect 1346 1526 1349 1596
rect 1354 1533 1365 1536
rect 1322 1513 1325 1526
rect 1338 1523 1349 1526
rect 1250 1373 1253 1423
rect 1258 1393 1261 1416
rect 1218 1353 1229 1356
rect 1218 1343 1221 1353
rect 1210 1313 1213 1326
rect 1202 1303 1213 1306
rect 1130 1213 1133 1226
rect 1066 1183 1069 1206
rect 1114 1203 1125 1206
rect 1146 1203 1149 1246
rect 1174 1243 1181 1246
rect 1170 1213 1173 1226
rect 1178 1196 1181 1243
rect 1186 1236 1189 1256
rect 1186 1233 1193 1236
rect 1174 1193 1181 1196
rect 1050 1003 1053 1136
rect 1058 1123 1061 1156
rect 1066 1033 1069 1176
rect 1058 1013 1061 1026
rect 1074 1013 1077 1136
rect 1090 1133 1093 1186
rect 1082 1113 1085 1126
rect 1098 1096 1101 1126
rect 1090 1093 1101 1096
rect 1090 1036 1093 1093
rect 1090 1033 1101 1036
rect 1098 1013 1101 1033
rect 1106 1006 1109 1186
rect 1114 1113 1117 1126
rect 1090 1003 1109 1006
rect 930 713 949 716
rect 930 593 933 616
rect 938 586 941 696
rect 946 613 949 713
rect 954 603 957 756
rect 962 723 965 836
rect 970 813 973 826
rect 970 733 973 746
rect 978 716 981 826
rect 986 723 989 816
rect 1010 813 1021 816
rect 1010 793 1013 806
rect 1018 746 1021 766
rect 1010 743 1021 746
rect 962 696 965 716
rect 978 713 989 716
rect 962 693 973 696
rect 970 636 973 693
rect 962 633 973 636
rect 898 583 925 586
rect 930 583 941 586
rect 842 443 845 536
rect 850 503 853 526
rect 858 463 861 536
rect 866 503 869 583
rect 874 513 877 566
rect 890 473 893 526
rect 898 493 901 526
rect 826 376 829 406
rect 842 403 845 426
rect 866 423 877 426
rect 898 423 901 436
rect 782 373 789 376
rect 786 353 789 373
rect 794 373 829 376
rect 746 213 749 226
rect 714 183 717 206
rect 722 193 725 206
rect 738 203 749 206
rect 706 123 709 136
rect 714 133 717 156
rect 746 153 749 203
rect 730 133 733 146
rect 762 143 765 206
rect 794 163 797 373
rect 850 366 853 416
rect 834 363 853 366
rect 834 316 837 363
rect 842 323 845 346
rect 834 313 845 316
rect 858 313 861 416
rect 866 383 869 406
rect 874 333 877 406
rect 882 403 885 416
rect 906 413 909 506
rect 922 483 925 536
rect 930 533 933 583
rect 962 553 965 633
rect 978 593 981 616
rect 986 603 989 713
rect 1010 646 1013 743
rect 1026 723 1029 806
rect 1034 716 1037 816
rect 1042 813 1045 826
rect 1042 733 1045 766
rect 1026 713 1037 716
rect 1010 643 1021 646
rect 1002 603 1005 626
rect 1010 596 1013 606
rect 986 593 1013 596
rect 1018 573 1021 643
rect 1026 603 1029 713
rect 1034 613 1037 706
rect 1042 703 1045 716
rect 1050 696 1053 936
rect 1066 933 1077 936
rect 1090 916 1093 1003
rect 1082 913 1093 916
rect 1058 893 1061 906
rect 1082 846 1085 913
rect 1098 896 1101 946
rect 1114 933 1117 1006
rect 1122 933 1125 1136
rect 1106 913 1109 926
rect 1098 893 1109 896
rect 1082 843 1093 846
rect 1058 793 1061 806
rect 1066 763 1069 826
rect 1082 753 1085 806
rect 1058 723 1061 746
rect 1090 736 1093 843
rect 1082 733 1093 736
rect 1042 693 1053 696
rect 1042 603 1045 693
rect 1082 686 1085 733
rect 1098 723 1101 826
rect 1106 813 1109 893
rect 1130 836 1133 996
rect 1138 853 1141 1166
rect 1162 1013 1165 1136
rect 1174 1006 1177 1193
rect 1190 1186 1193 1233
rect 1186 1183 1193 1186
rect 1146 903 1149 1006
rect 1174 1003 1181 1006
rect 1178 983 1181 1003
rect 1154 933 1181 936
rect 1170 903 1173 916
rect 1186 903 1189 1183
rect 1210 1133 1213 1303
rect 1218 1193 1221 1336
rect 1234 1286 1237 1336
rect 1266 1323 1269 1416
rect 1298 1413 1301 1436
rect 1306 1433 1309 1446
rect 1234 1283 1245 1286
rect 1226 1176 1229 1276
rect 1234 1213 1237 1266
rect 1242 1243 1245 1283
rect 1242 1213 1245 1226
rect 1226 1173 1237 1176
rect 1202 1046 1205 1126
rect 1210 1103 1213 1116
rect 1234 1096 1237 1173
rect 1258 1143 1261 1246
rect 1282 1213 1285 1226
rect 1290 1166 1293 1236
rect 1282 1163 1293 1166
rect 1194 1043 1205 1046
rect 1226 1093 1237 1096
rect 1194 1003 1197 1043
rect 1194 923 1197 936
rect 1202 923 1205 1016
rect 1226 973 1229 1093
rect 1282 1086 1285 1163
rect 1282 1083 1293 1086
rect 1298 1083 1301 1406
rect 1306 1123 1309 1426
rect 1314 1253 1317 1396
rect 1322 1333 1325 1486
rect 1354 1436 1357 1526
rect 1338 1433 1357 1436
rect 1330 1413 1333 1426
rect 1346 1413 1349 1426
rect 1362 1423 1365 1456
rect 1370 1443 1373 1616
rect 1378 1523 1381 1616
rect 1390 1613 1397 1616
rect 1390 1536 1393 1613
rect 1402 1576 1405 1606
rect 1410 1586 1413 1636
rect 1418 1623 1429 1626
rect 1418 1613 1445 1616
rect 1450 1603 1453 1636
rect 1458 1596 1461 1676
rect 1442 1593 1461 1596
rect 1410 1583 1421 1586
rect 1402 1573 1413 1576
rect 1386 1533 1393 1536
rect 1402 1533 1405 1566
rect 1386 1403 1389 1533
rect 1394 1513 1397 1526
rect 1402 1493 1405 1526
rect 1402 1413 1405 1426
rect 1410 1423 1413 1573
rect 1418 1533 1421 1583
rect 1418 1433 1421 1526
rect 1426 1433 1429 1536
rect 1434 1533 1437 1546
rect 1434 1513 1437 1526
rect 1442 1496 1445 1593
rect 1466 1536 1469 1656
rect 1438 1493 1445 1496
rect 1450 1533 1469 1536
rect 1438 1426 1441 1493
rect 1450 1443 1453 1533
rect 1458 1523 1469 1526
rect 1426 1423 1441 1426
rect 1370 1333 1373 1346
rect 1378 1333 1381 1356
rect 1402 1326 1405 1336
rect 1322 1166 1325 1326
rect 1318 1163 1325 1166
rect 1226 933 1229 946
rect 1234 933 1237 1026
rect 1242 963 1245 1036
rect 1250 1013 1261 1016
rect 1250 966 1253 1006
rect 1266 1003 1269 1026
rect 1274 966 1277 1066
rect 1290 1033 1293 1083
rect 1282 1003 1285 1016
rect 1298 1003 1301 1026
rect 1306 1013 1309 1106
rect 1318 1086 1321 1163
rect 1318 1083 1325 1086
rect 1322 1063 1325 1083
rect 1306 996 1309 1006
rect 1314 1003 1317 1056
rect 1330 1036 1333 1226
rect 1338 1146 1341 1316
rect 1386 1313 1389 1326
rect 1394 1323 1405 1326
rect 1410 1323 1413 1336
rect 1394 1306 1397 1323
rect 1418 1316 1421 1406
rect 1402 1313 1421 1316
rect 1394 1303 1405 1306
rect 1346 1213 1349 1236
rect 1346 1163 1349 1206
rect 1378 1153 1381 1186
rect 1394 1153 1397 1206
rect 1402 1203 1405 1303
rect 1426 1233 1429 1423
rect 1434 1333 1437 1416
rect 1442 1343 1445 1406
rect 1450 1336 1453 1416
rect 1458 1393 1461 1406
rect 1466 1403 1469 1416
rect 1458 1343 1461 1356
rect 1450 1333 1461 1336
rect 1426 1213 1429 1226
rect 1434 1213 1437 1306
rect 1442 1236 1445 1326
rect 1442 1233 1461 1236
rect 1458 1213 1461 1226
rect 1466 1223 1469 1346
rect 1474 1206 1477 1686
rect 1498 1676 1501 1716
rect 1498 1673 1517 1676
rect 1482 1603 1485 1616
rect 1490 1593 1493 1626
rect 1498 1583 1501 1666
rect 1506 1603 1509 1636
rect 1514 1623 1517 1673
rect 1522 1656 1525 1756
rect 1530 1713 1533 1726
rect 1522 1653 1533 1656
rect 1522 1633 1525 1646
rect 1482 1533 1501 1536
rect 1482 1513 1485 1526
rect 1490 1423 1493 1526
rect 1498 1493 1501 1533
rect 1506 1526 1509 1546
rect 1514 1543 1517 1616
rect 1522 1533 1525 1626
rect 1506 1523 1525 1526
rect 1514 1513 1525 1516
rect 1482 1373 1485 1416
rect 1490 1333 1493 1406
rect 1498 1393 1501 1416
rect 1482 1313 1485 1326
rect 1498 1316 1501 1376
rect 1514 1373 1517 1513
rect 1530 1423 1533 1653
rect 1538 1613 1541 1813
rect 1546 1673 1549 1736
rect 1554 1683 1557 1776
rect 1578 1746 1581 1843
rect 1602 1836 1605 1926
rect 1610 1923 1621 1926
rect 1610 1913 1613 1923
rect 1634 1913 1637 1926
rect 1642 1923 1653 1926
rect 1658 1906 1661 1926
rect 1654 1903 1661 1906
rect 1654 1836 1657 1903
rect 1602 1833 1613 1836
rect 1654 1833 1661 1836
rect 1570 1743 1581 1746
rect 1570 1686 1573 1743
rect 1570 1683 1581 1686
rect 1578 1663 1581 1683
rect 1546 1596 1549 1636
rect 1554 1623 1557 1656
rect 1554 1613 1565 1616
rect 1586 1613 1589 1736
rect 1594 1643 1597 1826
rect 1610 1776 1613 1833
rect 1642 1813 1645 1826
rect 1658 1813 1661 1833
rect 1666 1813 1669 1926
rect 1682 1906 1685 1916
rect 1690 1913 1693 1926
rect 1698 1906 1701 1996
rect 1710 1906 1713 2013
rect 1722 1943 1725 2006
rect 1738 1946 1741 2006
rect 1754 1966 1757 2093
rect 1778 2046 1781 2116
rect 1794 2103 1797 2216
rect 1802 2213 1805 2293
rect 1814 2236 1817 2303
rect 1810 2233 1817 2236
rect 1810 2213 1813 2233
rect 1826 2216 1829 2316
rect 1858 2246 1861 2326
rect 1882 2323 1885 2416
rect 1890 2323 1893 2423
rect 1922 2413 1925 2536
rect 1930 2423 1933 2526
rect 1946 2486 1949 2536
rect 1938 2483 1949 2486
rect 1938 2423 1941 2483
rect 1946 2423 1957 2426
rect 1962 2423 1965 2446
rect 1906 2356 1909 2406
rect 1922 2403 1941 2406
rect 1938 2393 1941 2403
rect 1898 2353 1909 2356
rect 1898 2323 1901 2353
rect 1906 2343 1933 2346
rect 1906 2333 1909 2343
rect 1914 2323 1917 2336
rect 1930 2333 1933 2343
rect 1946 2336 1949 2423
rect 1970 2416 1973 2526
rect 1978 2443 1981 2526
rect 2002 2433 2005 2543
rect 2010 2526 2013 2536
rect 2018 2533 2021 2543
rect 2026 2533 2037 2536
rect 2010 2523 2037 2526
rect 1954 2413 1973 2416
rect 1954 2346 1957 2413
rect 1962 2356 1965 2406
rect 1986 2393 1989 2406
rect 1994 2403 1997 2426
rect 2010 2406 2013 2456
rect 2018 2423 2021 2436
rect 2034 2416 2037 2516
rect 2042 2423 2045 2446
rect 2026 2413 2037 2416
rect 2050 2413 2069 2416
rect 2010 2403 2045 2406
rect 1962 2353 1973 2356
rect 1954 2343 1965 2346
rect 1946 2333 1957 2336
rect 1930 2323 1949 2326
rect 1954 2323 1957 2333
rect 1946 2316 1949 2323
rect 1850 2243 1861 2246
rect 1826 2213 1837 2216
rect 1802 2193 1805 2206
rect 1818 2203 1829 2206
rect 1834 2193 1837 2213
rect 1802 2163 1829 2166
rect 1802 2133 1805 2163
rect 1810 2113 1813 2156
rect 1826 2153 1829 2163
rect 1818 2133 1829 2136
rect 1818 2113 1821 2126
rect 1826 2113 1829 2133
rect 1834 2123 1837 2136
rect 1842 2133 1845 2226
rect 1850 2153 1853 2243
rect 1858 2203 1861 2236
rect 1866 2193 1869 2206
rect 1874 2173 1877 2226
rect 1882 2116 1885 2226
rect 1906 2213 1909 2226
rect 1922 2223 1925 2286
rect 1890 2183 1893 2206
rect 1890 2133 1893 2156
rect 1770 2043 1781 2046
rect 1754 1963 1761 1966
rect 1738 1943 1749 1946
rect 1730 1933 1741 1936
rect 1682 1903 1701 1906
rect 1706 1903 1713 1906
rect 1682 1836 1685 1903
rect 1706 1886 1709 1903
rect 1674 1833 1685 1836
rect 1698 1883 1709 1886
rect 1634 1793 1637 1806
rect 1602 1773 1613 1776
rect 1602 1753 1605 1773
rect 1546 1593 1553 1596
rect 1538 1523 1541 1586
rect 1538 1503 1541 1516
rect 1550 1496 1553 1593
rect 1562 1533 1565 1606
rect 1610 1603 1613 1726
rect 1642 1713 1645 1736
rect 1650 1733 1653 1806
rect 1674 1803 1677 1833
rect 1682 1803 1685 1826
rect 1698 1746 1701 1883
rect 1722 1876 1725 1926
rect 1730 1913 1733 1926
rect 1746 1903 1749 1943
rect 1714 1873 1725 1876
rect 1706 1793 1709 1806
rect 1714 1793 1717 1873
rect 1730 1813 1733 1826
rect 1746 1793 1749 1806
rect 1758 1756 1761 1963
rect 1758 1753 1765 1756
rect 1770 1753 1773 2043
rect 1778 2023 1781 2036
rect 1786 1933 1789 2016
rect 1778 1803 1781 1916
rect 1794 1896 1797 2066
rect 1818 2013 1837 2016
rect 1802 1983 1805 2006
rect 1810 2003 1821 2006
rect 1810 1923 1813 2003
rect 1786 1893 1797 1896
rect 1786 1793 1789 1893
rect 1794 1803 1797 1886
rect 1818 1813 1821 1946
rect 1826 1933 1829 2006
rect 1834 1823 1837 2013
rect 1842 1903 1845 1976
rect 1850 1873 1853 2116
rect 1882 2113 1893 2116
rect 1874 2103 1885 2106
rect 1866 2003 1869 2016
rect 1874 1996 1877 2066
rect 1906 2063 1909 2186
rect 1922 2096 1925 2186
rect 1938 2166 1941 2316
rect 1946 2313 1957 2316
rect 1962 2303 1965 2343
rect 1970 2313 1973 2353
rect 2018 2343 2021 2386
rect 2050 2383 2053 2406
rect 2074 2403 2085 2406
rect 2090 2403 2093 2536
rect 2098 2533 2101 2546
rect 2098 2423 2101 2436
rect 2098 2386 2101 2416
rect 2130 2413 2133 2526
rect 2162 2433 2165 2536
rect 2170 2483 2173 2536
rect 2178 2413 2181 2526
rect 2114 2403 2125 2406
rect 2106 2393 2117 2396
rect 2098 2383 2109 2386
rect 2114 2383 2117 2393
rect 2026 2333 2029 2376
rect 2042 2333 2053 2336
rect 1978 2313 1981 2326
rect 1986 2323 2005 2326
rect 1986 2303 1989 2323
rect 1946 2203 1949 2256
rect 1970 2213 1973 2226
rect 1930 2163 1941 2166
rect 1930 2133 1933 2163
rect 1978 2096 1981 2186
rect 1994 2176 1997 2316
rect 2050 2296 2053 2326
rect 2082 2323 2101 2326
rect 2074 2313 2085 2316
rect 2106 2303 2109 2383
rect 2042 2293 2053 2296
rect 2042 2246 2045 2293
rect 2042 2243 2053 2246
rect 1986 2173 1997 2176
rect 2002 2173 2005 2206
rect 2050 2203 2053 2243
rect 2058 2186 2061 2216
rect 2066 2203 2069 2286
rect 2098 2213 2101 2226
rect 2122 2203 2125 2316
rect 2170 2186 2173 2366
rect 2186 2346 2189 2416
rect 2194 2363 2197 2406
rect 2242 2373 2245 2406
rect 2250 2393 2253 2546
rect 2274 2543 2301 2546
rect 2274 2536 2277 2543
rect 2266 2533 2277 2536
rect 2282 2533 2293 2536
rect 2298 2533 2301 2543
rect 2266 2413 2269 2533
rect 2274 2523 2293 2526
rect 2298 2513 2301 2526
rect 2186 2343 2197 2346
rect 2202 2343 2205 2356
rect 2194 2336 2197 2343
rect 2178 2313 2181 2326
rect 2034 2183 2061 2186
rect 2090 2183 2101 2186
rect 2170 2183 2181 2186
rect 1986 2133 1989 2173
rect 1922 2093 1933 2096
rect 1882 2013 1885 2026
rect 1890 2003 1893 2016
rect 1874 1993 1893 1996
rect 1834 1756 1837 1806
rect 1818 1753 1837 1756
rect 1842 1753 1845 1826
rect 1850 1823 1853 1836
rect 1858 1833 1861 1946
rect 1882 1933 1885 1956
rect 1866 1826 1869 1926
rect 1874 1883 1877 1916
rect 1882 1903 1885 1916
rect 1890 1893 1893 1993
rect 1906 1973 1909 2016
rect 1914 1953 1917 2036
rect 1922 1946 1925 2026
rect 1930 1963 1933 2093
rect 1962 2093 1981 2096
rect 1962 2006 1965 2093
rect 1938 1953 1941 2006
rect 1962 2003 1981 2006
rect 1978 1983 1981 2003
rect 1986 1953 1989 2126
rect 2010 2013 2013 2026
rect 2034 2003 2037 2183
rect 2042 2133 2045 2176
rect 2042 2096 2045 2126
rect 2042 2093 2049 2096
rect 2046 2026 2049 2093
rect 2042 2023 2049 2026
rect 1914 1943 1925 1946
rect 1858 1823 1869 1826
rect 1858 1813 1861 1823
rect 1698 1743 1709 1746
rect 1674 1713 1677 1726
rect 1618 1613 1621 1626
rect 1634 1613 1637 1676
rect 1650 1623 1653 1646
rect 1570 1496 1573 1516
rect 1546 1493 1553 1496
rect 1562 1493 1573 1496
rect 1506 1323 1509 1356
rect 1514 1316 1517 1326
rect 1498 1313 1517 1316
rect 1514 1293 1517 1313
rect 1522 1276 1525 1416
rect 1546 1406 1549 1493
rect 1562 1446 1565 1493
rect 1562 1443 1573 1446
rect 1530 1403 1549 1406
rect 1530 1333 1533 1403
rect 1554 1396 1557 1426
rect 1546 1393 1557 1396
rect 1562 1393 1565 1416
rect 1538 1326 1541 1376
rect 1514 1273 1525 1276
rect 1534 1323 1541 1326
rect 1338 1143 1349 1146
rect 1346 1076 1349 1143
rect 1338 1073 1349 1076
rect 1338 1053 1341 1073
rect 1322 996 1325 1036
rect 1330 1033 1341 1036
rect 1282 993 1309 996
rect 1314 993 1325 996
rect 1250 963 1261 966
rect 1258 933 1261 963
rect 1266 963 1277 966
rect 1218 893 1221 926
rect 1234 906 1237 926
rect 1242 913 1245 926
rect 1122 833 1133 836
rect 1122 813 1125 833
rect 1138 813 1141 826
rect 1106 693 1109 736
rect 1122 733 1125 806
rect 1082 683 1093 686
rect 1066 613 1069 626
rect 1090 563 1093 683
rect 1130 676 1133 776
rect 1138 723 1141 756
rect 1170 753 1173 826
rect 1178 773 1181 806
rect 1226 773 1229 906
rect 1234 903 1245 906
rect 1234 813 1237 896
rect 1266 893 1269 963
rect 1274 943 1277 956
rect 1282 926 1285 966
rect 1278 923 1285 926
rect 1278 846 1281 923
rect 1290 863 1293 946
rect 1278 843 1285 846
rect 1258 813 1261 826
rect 1282 786 1285 843
rect 1290 803 1293 856
rect 1298 833 1301 986
rect 1314 953 1317 993
rect 1306 913 1309 926
rect 1322 893 1325 976
rect 1330 906 1333 1026
rect 1338 946 1341 1033
rect 1354 1013 1357 1036
rect 1370 1013 1373 1126
rect 1386 1093 1389 1136
rect 1458 1133 1461 1206
rect 1470 1203 1477 1206
rect 1470 1096 1473 1203
rect 1482 1106 1485 1236
rect 1490 1113 1493 1126
rect 1498 1113 1501 1226
rect 1514 1186 1517 1273
rect 1534 1266 1537 1323
rect 1546 1283 1549 1393
rect 1570 1336 1573 1443
rect 1578 1433 1581 1556
rect 1594 1496 1597 1586
rect 1618 1566 1621 1606
rect 1666 1603 1669 1696
rect 1698 1643 1701 1736
rect 1706 1673 1709 1743
rect 1730 1636 1733 1726
rect 1738 1693 1741 1726
rect 1754 1723 1757 1736
rect 1762 1713 1765 1753
rect 1786 1716 1789 1726
rect 1778 1713 1789 1716
rect 1794 1713 1797 1726
rect 1778 1683 1781 1713
rect 1674 1613 1677 1636
rect 1722 1633 1733 1636
rect 1610 1563 1621 1566
rect 1634 1563 1637 1586
rect 1610 1506 1613 1563
rect 1650 1556 1653 1586
rect 1650 1553 1661 1556
rect 1586 1493 1597 1496
rect 1602 1503 1613 1506
rect 1586 1413 1589 1493
rect 1602 1486 1605 1503
rect 1626 1496 1629 1526
rect 1658 1523 1661 1553
rect 1594 1483 1605 1486
rect 1610 1493 1629 1496
rect 1666 1493 1669 1596
rect 1674 1553 1677 1606
rect 1722 1583 1725 1633
rect 1730 1603 1733 1626
rect 1762 1613 1765 1626
rect 1778 1603 1781 1616
rect 1786 1603 1789 1706
rect 1810 1703 1813 1736
rect 1810 1613 1813 1636
rect 1818 1613 1821 1753
rect 1842 1703 1845 1726
rect 1834 1603 1837 1636
rect 1842 1596 1845 1696
rect 1866 1636 1869 1736
rect 1874 1733 1877 1876
rect 1898 1833 1901 1916
rect 1906 1913 1909 1936
rect 1914 1923 1917 1943
rect 1922 1923 1925 1936
rect 1906 1833 1909 1906
rect 1890 1813 1893 1826
rect 1898 1813 1901 1826
rect 1874 1693 1877 1726
rect 1898 1713 1901 1726
rect 1866 1633 1877 1636
rect 1866 1613 1869 1626
rect 1874 1613 1877 1633
rect 1834 1593 1845 1596
rect 1594 1403 1597 1483
rect 1602 1396 1605 1406
rect 1578 1393 1605 1396
rect 1602 1346 1605 1393
rect 1610 1356 1613 1493
rect 1642 1426 1645 1446
rect 1626 1413 1629 1426
rect 1638 1423 1645 1426
rect 1610 1353 1629 1356
rect 1602 1343 1613 1346
rect 1530 1263 1537 1266
rect 1530 1193 1533 1263
rect 1554 1216 1557 1326
rect 1562 1223 1565 1336
rect 1570 1333 1581 1336
rect 1570 1313 1573 1326
rect 1578 1276 1581 1333
rect 1586 1313 1589 1336
rect 1594 1323 1597 1336
rect 1602 1293 1605 1336
rect 1610 1323 1613 1343
rect 1618 1333 1621 1346
rect 1578 1273 1589 1276
rect 1538 1213 1557 1216
rect 1514 1183 1525 1186
rect 1506 1113 1509 1156
rect 1482 1103 1509 1106
rect 1522 1103 1525 1183
rect 1538 1103 1541 1213
rect 1586 1206 1589 1273
rect 1546 1113 1549 1206
rect 1554 1203 1589 1206
rect 1554 1113 1557 1203
rect 1610 1196 1613 1286
rect 1618 1203 1621 1326
rect 1562 1133 1565 1196
rect 1610 1193 1621 1196
rect 1626 1193 1629 1353
rect 1638 1346 1641 1423
rect 1638 1343 1645 1346
rect 1642 1326 1645 1343
rect 1650 1333 1653 1416
rect 1642 1323 1653 1326
rect 1658 1323 1661 1336
rect 1634 1303 1637 1316
rect 1650 1256 1653 1323
rect 1666 1313 1669 1326
rect 1674 1323 1677 1336
rect 1646 1253 1653 1256
rect 1610 1133 1613 1156
rect 1618 1133 1621 1193
rect 1634 1153 1637 1216
rect 1646 1176 1649 1253
rect 1682 1236 1685 1526
rect 1714 1513 1717 1536
rect 1722 1533 1725 1566
rect 1746 1513 1749 1526
rect 1770 1463 1773 1536
rect 1722 1296 1725 1366
rect 1754 1333 1757 1346
rect 1730 1313 1733 1326
rect 1770 1313 1773 1326
rect 1778 1323 1781 1546
rect 1802 1503 1805 1526
rect 1826 1523 1829 1536
rect 1834 1533 1837 1593
rect 1874 1553 1877 1586
rect 1858 1513 1861 1526
rect 1882 1473 1885 1536
rect 1890 1456 1893 1636
rect 1898 1543 1901 1646
rect 1882 1453 1893 1456
rect 1794 1363 1813 1366
rect 1794 1333 1797 1363
rect 1722 1293 1741 1296
rect 1674 1233 1685 1236
rect 1674 1176 1677 1233
rect 1690 1213 1693 1226
rect 1730 1213 1733 1226
rect 1646 1173 1653 1176
rect 1674 1173 1709 1176
rect 1650 1153 1653 1173
rect 1470 1093 1477 1096
rect 1386 1003 1389 1036
rect 1394 1003 1397 1086
rect 1474 1013 1477 1093
rect 1482 1013 1485 1036
rect 1410 983 1421 986
rect 1338 943 1349 946
rect 1338 913 1341 936
rect 1346 923 1349 943
rect 1354 933 1357 956
rect 1370 933 1373 946
rect 1330 903 1349 906
rect 1354 903 1357 916
rect 1386 883 1389 926
rect 1338 803 1341 826
rect 1258 783 1285 786
rect 1126 673 1133 676
rect 1126 626 1129 673
rect 1146 666 1149 736
rect 1194 733 1197 746
rect 1202 733 1205 756
rect 1250 733 1253 766
rect 1258 733 1261 783
rect 1298 753 1301 786
rect 1138 663 1149 666
rect 1098 593 1101 606
rect 930 493 933 526
rect 946 496 949 516
rect 942 493 949 496
rect 898 366 901 406
rect 914 403 917 446
rect 922 413 925 426
rect 930 403 933 466
rect 890 363 901 366
rect 942 366 945 493
rect 942 363 949 366
rect 882 316 885 356
rect 890 343 893 363
rect 890 323 893 336
rect 898 333 901 356
rect 898 316 901 326
rect 882 313 901 316
rect 810 193 813 216
rect 778 123 781 146
rect 826 113 829 126
rect 842 123 845 313
rect 946 296 949 363
rect 938 293 949 296
rect 858 213 861 226
rect 874 216 877 236
rect 938 226 941 293
rect 874 213 893 216
rect 890 193 893 206
rect 898 203 901 226
rect 938 223 949 226
rect 850 126 853 156
rect 858 133 861 146
rect 874 133 877 166
rect 906 133 909 206
rect 930 166 933 206
rect 922 163 933 166
rect 850 123 861 126
rect 922 123 925 163
rect 858 113 861 123
rect 946 113 949 223
rect 954 213 957 526
rect 978 443 981 536
rect 1002 493 1005 526
rect 962 403 965 416
rect 962 293 965 356
rect 970 316 973 416
rect 978 333 981 426
rect 994 413 997 436
rect 986 383 989 406
rect 1002 336 1005 416
rect 1010 413 1013 526
rect 1034 523 1037 536
rect 1002 333 1013 336
rect 970 313 981 316
rect 978 236 981 313
rect 962 223 965 236
rect 970 233 981 236
rect 970 196 973 233
rect 978 203 981 216
rect 970 193 981 196
rect 970 123 973 136
rect 690 103 701 106
rect 978 103 981 193
rect 986 153 989 216
rect 994 183 997 206
rect 1002 203 1005 333
rect 1010 193 1013 216
rect 1018 213 1021 416
rect 1026 403 1029 506
rect 1042 423 1045 536
rect 1090 533 1093 556
rect 1106 543 1109 606
rect 1114 536 1117 626
rect 1126 623 1133 626
rect 1130 603 1133 623
rect 1138 596 1141 663
rect 1146 603 1149 616
rect 1138 593 1149 596
rect 1106 533 1117 536
rect 1066 473 1069 526
rect 1098 513 1101 526
rect 1106 496 1109 533
rect 1098 493 1109 496
rect 1082 423 1085 446
rect 1098 426 1101 493
rect 1114 456 1117 526
rect 1122 503 1125 536
rect 1130 503 1133 516
rect 1138 456 1141 546
rect 1146 503 1149 593
rect 1154 533 1157 616
rect 1154 513 1157 526
rect 1114 453 1125 456
rect 1098 423 1109 426
rect 1114 423 1117 436
rect 1026 323 1029 376
rect 1034 306 1037 326
rect 1030 303 1037 306
rect 1030 196 1033 303
rect 1042 233 1045 326
rect 1042 203 1045 216
rect 1030 193 1037 196
rect 1026 133 1029 166
rect 994 113 997 126
rect 666 93 677 96
rect 674 -96 677 93
rect 698 16 701 103
rect 1034 93 1037 193
rect 1050 183 1053 386
rect 1098 383 1101 406
rect 1106 373 1109 423
rect 1122 416 1125 453
rect 1130 453 1141 456
rect 1162 453 1165 606
rect 1170 493 1173 616
rect 1178 523 1181 606
rect 1186 603 1189 626
rect 1186 533 1189 596
rect 1130 423 1133 453
rect 1186 423 1189 436
rect 1122 413 1141 416
rect 1114 403 1125 406
rect 1162 403 1165 416
rect 1058 253 1061 366
rect 1114 333 1117 346
rect 1122 333 1125 403
rect 1058 153 1061 216
rect 1066 203 1069 266
rect 1082 213 1085 326
rect 1090 313 1093 326
rect 1130 323 1133 396
rect 1170 383 1173 406
rect 1178 393 1181 406
rect 1138 313 1141 336
rect 1162 213 1165 326
rect 1194 323 1197 646
rect 1202 403 1205 566
rect 1210 556 1213 616
rect 1226 593 1229 726
rect 1234 603 1237 626
rect 1210 553 1221 556
rect 1210 523 1213 546
rect 1210 403 1213 516
rect 1218 513 1221 553
rect 1242 543 1245 616
rect 1258 596 1261 616
rect 1250 593 1261 596
rect 1250 536 1253 593
rect 1266 563 1269 626
rect 1282 623 1285 726
rect 1274 536 1277 596
rect 1298 536 1301 706
rect 1306 623 1309 736
rect 1314 713 1317 786
rect 1346 763 1349 806
rect 1394 803 1397 926
rect 1410 853 1413 906
rect 1418 846 1421 983
rect 1442 963 1445 1006
rect 1450 993 1453 1006
rect 1426 923 1429 936
rect 1450 916 1453 926
rect 1442 913 1453 916
rect 1410 843 1421 846
rect 1402 783 1405 816
rect 1410 786 1413 843
rect 1418 793 1421 816
rect 1426 803 1429 896
rect 1450 873 1453 913
rect 1474 836 1477 956
rect 1482 933 1485 986
rect 1498 953 1501 1036
rect 1506 1013 1509 1103
rect 1530 1013 1533 1026
rect 1506 993 1509 1006
rect 1554 1003 1557 1016
rect 1562 1003 1565 1126
rect 1586 1013 1589 1026
rect 1610 1003 1613 1016
rect 1482 893 1485 926
rect 1506 913 1509 926
rect 1530 843 1533 936
rect 1538 933 1541 986
rect 1618 983 1621 1126
rect 1642 1066 1645 1126
rect 1666 1123 1669 1136
rect 1682 1133 1685 1146
rect 1634 1063 1645 1066
rect 1634 1013 1637 1063
rect 1642 1013 1645 1036
rect 1642 933 1645 986
rect 1666 953 1669 1026
rect 1674 1003 1677 1086
rect 1706 1083 1709 1173
rect 1714 1126 1717 1206
rect 1738 1183 1741 1293
rect 1786 1256 1789 1326
rect 1802 1323 1805 1336
rect 1810 1323 1813 1363
rect 1778 1253 1789 1256
rect 1730 1143 1733 1166
rect 1714 1123 1721 1126
rect 1718 1036 1721 1123
rect 1730 1113 1733 1126
rect 1746 1053 1749 1216
rect 1770 1196 1773 1206
rect 1778 1203 1781 1253
rect 1786 1196 1789 1216
rect 1770 1193 1789 1196
rect 1754 1123 1765 1126
rect 1718 1033 1741 1036
rect 1698 1013 1701 1026
rect 1722 993 1725 1006
rect 1738 1003 1741 1033
rect 1562 893 1565 926
rect 1474 833 1493 836
rect 1474 823 1485 826
rect 1482 803 1485 816
rect 1490 793 1493 833
rect 1506 823 1509 836
rect 1506 803 1509 816
rect 1410 783 1421 786
rect 1338 666 1341 726
rect 1362 706 1365 756
rect 1370 713 1373 736
rect 1418 733 1421 783
rect 1426 733 1429 776
rect 1514 753 1517 826
rect 1522 813 1533 816
rect 1538 813 1541 826
rect 1490 733 1493 746
rect 1514 733 1517 746
rect 1362 703 1373 706
rect 1394 703 1397 726
rect 1402 713 1405 726
rect 1338 663 1357 666
rect 1354 603 1357 663
rect 1362 613 1365 626
rect 1370 603 1373 703
rect 1450 623 1453 636
rect 1418 593 1421 606
rect 1426 603 1429 616
rect 1450 606 1453 616
rect 1474 613 1477 726
rect 1506 713 1509 726
rect 1442 593 1445 606
rect 1450 603 1477 606
rect 1490 603 1493 626
rect 1498 613 1501 646
rect 1506 623 1509 636
rect 1514 623 1517 706
rect 1522 646 1525 806
rect 1530 683 1533 813
rect 1538 733 1541 796
rect 1546 766 1549 886
rect 1586 883 1589 926
rect 1594 873 1597 926
rect 1554 813 1557 826
rect 1562 813 1565 826
rect 1570 796 1573 836
rect 1578 803 1581 816
rect 1586 806 1589 826
rect 1594 813 1597 826
rect 1586 803 1605 806
rect 1610 803 1613 816
rect 1618 813 1621 926
rect 1642 863 1645 926
rect 1650 913 1653 936
rect 1698 933 1701 956
rect 1706 933 1709 946
rect 1570 793 1581 796
rect 1546 763 1557 766
rect 1538 713 1541 726
rect 1546 703 1549 756
rect 1554 733 1557 763
rect 1522 643 1533 646
rect 1522 593 1525 606
rect 1530 603 1533 643
rect 1538 613 1541 666
rect 1546 613 1549 626
rect 1554 606 1557 716
rect 1562 663 1565 746
rect 1570 706 1573 736
rect 1578 723 1581 793
rect 1602 763 1605 803
rect 1570 703 1577 706
rect 1562 623 1565 656
rect 1574 636 1577 703
rect 1570 633 1577 636
rect 1570 616 1573 633
rect 1586 623 1589 736
rect 1546 603 1557 606
rect 1562 613 1573 616
rect 1562 603 1565 613
rect 1586 603 1589 616
rect 1594 603 1597 626
rect 1602 613 1605 726
rect 1610 636 1613 716
rect 1610 633 1621 636
rect 1610 606 1613 616
rect 1602 603 1613 606
rect 1618 606 1621 633
rect 1626 613 1629 636
rect 1634 613 1637 806
rect 1642 803 1645 816
rect 1658 766 1661 826
rect 1666 773 1669 926
rect 1706 896 1709 916
rect 1730 913 1733 926
rect 1706 893 1717 896
rect 1698 813 1701 826
rect 1658 763 1669 766
rect 1650 683 1661 686
rect 1650 613 1653 646
rect 1658 613 1661 683
rect 1666 653 1669 763
rect 1674 676 1677 786
rect 1714 783 1717 893
rect 1722 813 1725 896
rect 1746 813 1749 866
rect 1754 813 1757 936
rect 1762 833 1765 1123
rect 1770 1113 1773 1126
rect 1770 863 1773 1056
rect 1778 996 1781 1156
rect 1794 1153 1797 1266
rect 1818 1263 1821 1336
rect 1826 1323 1829 1336
rect 1858 1333 1861 1406
rect 1882 1403 1885 1453
rect 1890 1403 1893 1416
rect 1898 1413 1901 1536
rect 1906 1453 1909 1726
rect 1922 1653 1925 1836
rect 1930 1733 1933 1826
rect 1938 1666 1941 1826
rect 1946 1803 1949 1926
rect 1970 1813 1973 1926
rect 1978 1823 1981 1936
rect 2026 1933 2029 1986
rect 2042 1936 2045 2023
rect 2034 1933 2045 1936
rect 2034 1926 2037 1933
rect 2002 1903 2005 1926
rect 2026 1923 2037 1926
rect 2026 1896 2029 1923
rect 2034 1903 2037 1916
rect 1994 1746 1997 1806
rect 1986 1743 1997 1746
rect 1962 1673 1965 1726
rect 1938 1663 1965 1666
rect 1914 1593 1917 1606
rect 1914 1503 1917 1556
rect 1922 1523 1925 1586
rect 1930 1563 1933 1606
rect 1954 1583 1957 1616
rect 1938 1556 1941 1576
rect 1962 1573 1965 1663
rect 1930 1553 1941 1556
rect 1970 1553 1973 1656
rect 1986 1653 1989 1743
rect 1930 1533 1933 1553
rect 1946 1496 1949 1526
rect 1938 1493 1949 1496
rect 1938 1436 1941 1493
rect 1938 1433 1949 1436
rect 1858 1306 1861 1326
rect 1866 1323 1869 1336
rect 1850 1303 1861 1306
rect 1850 1246 1853 1303
rect 1850 1243 1861 1246
rect 1802 1126 1805 1236
rect 1810 1213 1813 1226
rect 1834 1213 1837 1226
rect 1858 1213 1861 1243
rect 1874 1226 1877 1356
rect 1882 1343 1901 1346
rect 1882 1323 1885 1343
rect 1890 1313 1893 1336
rect 1898 1333 1901 1343
rect 1866 1223 1877 1226
rect 1810 1183 1813 1206
rect 1866 1163 1869 1223
rect 1874 1183 1877 1216
rect 1898 1213 1901 1326
rect 1906 1273 1909 1406
rect 1914 1353 1917 1416
rect 1946 1413 1949 1433
rect 1930 1333 1933 1346
rect 1954 1343 1957 1526
rect 1962 1496 1965 1516
rect 1962 1493 1969 1496
rect 1914 1313 1917 1326
rect 1954 1313 1957 1326
rect 1966 1306 1969 1493
rect 1978 1333 1981 1596
rect 1994 1546 1997 1736
rect 2002 1673 2005 1816
rect 2010 1803 2013 1886
rect 2018 1783 2021 1896
rect 2026 1893 2037 1896
rect 2042 1893 2045 1926
rect 2050 1903 2053 2006
rect 2034 1886 2037 1893
rect 2058 1886 2061 2016
rect 2074 1986 2077 2026
rect 2066 1983 2077 1986
rect 2066 1893 2069 1983
rect 2026 1803 2029 1886
rect 2034 1883 2045 1886
rect 2058 1883 2069 1886
rect 2074 1883 2077 1936
rect 2034 1813 2037 1826
rect 2042 1786 2045 1883
rect 2050 1796 2053 1836
rect 2058 1813 2061 1826
rect 2066 1803 2069 1883
rect 2082 1826 2085 1916
rect 2090 1863 2093 2183
rect 2146 2133 2149 2146
rect 2130 2056 2133 2126
rect 2146 2113 2149 2126
rect 2154 2096 2157 2126
rect 2146 2093 2157 2096
rect 2130 2053 2137 2056
rect 2122 2013 2125 2046
rect 2098 1923 2101 1936
rect 2106 1853 2109 2006
rect 2082 1823 2101 1826
rect 2106 1823 2109 1846
rect 2074 1803 2077 1816
rect 2050 1793 2069 1796
rect 2042 1783 2053 1786
rect 2050 1733 2053 1783
rect 2058 1733 2061 1786
rect 2066 1736 2069 1793
rect 2066 1733 2077 1736
rect 1986 1543 1997 1546
rect 1986 1383 1989 1543
rect 1994 1523 1997 1536
rect 2002 1533 2005 1656
rect 2010 1613 2013 1636
rect 2018 1613 2021 1726
rect 2026 1706 2029 1726
rect 2066 1723 2069 1733
rect 2026 1703 2033 1706
rect 2030 1636 2033 1703
rect 2026 1633 2033 1636
rect 2018 1593 2021 1606
rect 2026 1553 2029 1633
rect 2034 1556 2037 1616
rect 2058 1613 2061 1626
rect 2082 1586 2085 1806
rect 2090 1783 2093 1823
rect 2114 1813 2117 2006
rect 2134 1986 2137 2053
rect 2146 2046 2149 2093
rect 2146 2043 2157 2046
rect 2162 2043 2165 2136
rect 2130 1983 2137 1986
rect 2130 1963 2133 1983
rect 2146 1956 2149 2006
rect 2130 1953 2149 1956
rect 2154 1953 2157 2043
rect 2162 1983 2165 1996
rect 2170 1976 2173 2146
rect 2178 2133 2181 2183
rect 2186 2073 2189 2336
rect 2194 2333 2205 2336
rect 2234 2333 2237 2356
rect 2242 2343 2245 2366
rect 2210 2303 2213 2326
rect 2210 2213 2213 2246
rect 2218 2236 2221 2326
rect 2218 2233 2229 2236
rect 2194 2103 2197 2136
rect 2218 2133 2221 2216
rect 2226 2213 2229 2233
rect 2234 2216 2237 2316
rect 2242 2313 2245 2336
rect 2258 2323 2261 2336
rect 2282 2333 2285 2436
rect 2250 2223 2253 2246
rect 2234 2213 2253 2216
rect 2274 2213 2277 2326
rect 2298 2313 2301 2416
rect 2306 2393 2309 2536
rect 2314 2533 2317 2546
rect 2322 2533 2349 2536
rect 2378 2533 2381 2546
rect 2322 2526 2325 2533
rect 2314 2523 2325 2526
rect 2314 2433 2317 2523
rect 2322 2476 2325 2516
rect 2330 2496 2333 2526
rect 2338 2503 2341 2516
rect 2346 2513 2349 2533
rect 2330 2493 2349 2496
rect 2354 2493 2357 2526
rect 2362 2503 2365 2516
rect 2322 2473 2333 2476
rect 2314 2403 2317 2416
rect 2330 2396 2333 2473
rect 2346 2413 2349 2493
rect 2370 2423 2373 2526
rect 2402 2523 2405 2556
rect 2410 2513 2413 2536
rect 2418 2523 2429 2526
rect 2418 2503 2421 2523
rect 2330 2393 2341 2396
rect 2330 2346 2333 2393
rect 2370 2383 2373 2406
rect 2378 2393 2381 2406
rect 2426 2403 2429 2516
rect 2434 2493 2437 2536
rect 2450 2533 2453 2556
rect 2466 2533 2493 2536
rect 2442 2513 2445 2526
rect 2466 2523 2469 2533
rect 2474 2503 2477 2526
rect 2482 2513 2485 2526
rect 2490 2453 2493 2533
rect 2498 2446 2501 2546
rect 2506 2513 2509 2526
rect 2490 2443 2501 2446
rect 2322 2343 2333 2346
rect 2322 2323 2325 2343
rect 2338 2336 2341 2366
rect 2330 2333 2341 2336
rect 2346 2306 2349 2376
rect 2434 2363 2437 2416
rect 2474 2406 2477 2416
rect 2490 2413 2493 2443
rect 2498 2413 2501 2426
rect 2338 2303 2349 2306
rect 2354 2333 2373 2336
rect 2338 2246 2341 2303
rect 2322 2243 2341 2246
rect 2226 2193 2229 2206
rect 2234 2203 2245 2206
rect 2234 2116 2237 2203
rect 2210 2113 2237 2116
rect 2250 2113 2253 2213
rect 2258 2133 2261 2146
rect 2210 2093 2213 2113
rect 2282 2083 2285 2156
rect 2290 2113 2293 2186
rect 2306 2126 2309 2136
rect 2298 2123 2309 2126
rect 2186 2013 2189 2026
rect 2162 1973 2173 1976
rect 2122 1913 2125 1926
rect 2130 1906 2133 1953
rect 2146 1933 2149 1946
rect 2154 1916 2157 1936
rect 2162 1933 2165 1973
rect 2126 1903 2133 1906
rect 2138 1903 2141 1916
rect 2150 1913 2157 1916
rect 2126 1846 2129 1903
rect 2122 1843 2129 1846
rect 2098 1793 2101 1806
rect 2114 1766 2117 1806
rect 2106 1763 2117 1766
rect 2106 1723 2109 1763
rect 2122 1706 2125 1843
rect 2150 1836 2153 1913
rect 2150 1833 2157 1836
rect 2130 1816 2133 1826
rect 2130 1813 2149 1816
rect 2130 1803 2141 1806
rect 2130 1733 2133 1803
rect 2138 1783 2141 1796
rect 2130 1716 2133 1726
rect 2130 1713 2141 1716
rect 2146 1713 2149 1813
rect 2154 1773 2157 1833
rect 2162 1813 2165 1916
rect 2170 1823 2173 1966
rect 2210 1926 2213 1956
rect 2218 1933 2221 2006
rect 2226 2003 2229 2026
rect 2226 1933 2229 1956
rect 2210 1923 2221 1926
rect 2218 1913 2221 1923
rect 2226 1913 2229 1926
rect 2234 1923 2237 2016
rect 2242 2013 2253 2016
rect 2178 1816 2181 1896
rect 2242 1893 2245 2013
rect 2250 1983 2253 2006
rect 2258 1976 2261 2026
rect 2250 1973 2261 1976
rect 2250 1903 2253 1973
rect 2186 1823 2189 1836
rect 2170 1813 2189 1816
rect 2058 1583 2085 1586
rect 2034 1553 2053 1556
rect 1994 1323 1997 1506
rect 1962 1303 1969 1306
rect 1930 1213 1933 1226
rect 1810 1143 1829 1146
rect 1810 1133 1813 1143
rect 1818 1126 1821 1136
rect 1794 1113 1797 1126
rect 1802 1123 1821 1126
rect 1826 1123 1829 1143
rect 1818 1053 1821 1123
rect 1834 1033 1837 1156
rect 1882 1153 1885 1206
rect 1930 1193 1933 1206
rect 1938 1203 1941 1216
rect 1962 1213 1965 1303
rect 1842 1073 1845 1136
rect 1898 1133 1901 1186
rect 1850 1113 1853 1126
rect 1874 1113 1877 1126
rect 1786 1013 1789 1026
rect 1810 1013 1821 1016
rect 1826 1013 1829 1026
rect 1842 1013 1853 1016
rect 1778 993 1785 996
rect 1782 916 1785 993
rect 1834 976 1837 996
rect 1830 973 1837 976
rect 1778 913 1785 916
rect 1778 893 1781 913
rect 1722 766 1725 796
rect 1682 713 1685 766
rect 1714 763 1725 766
rect 1690 723 1693 736
rect 1714 686 1717 763
rect 1730 733 1733 746
rect 1714 683 1725 686
rect 1674 673 1685 676
rect 1618 603 1637 606
rect 1642 603 1653 606
rect 1658 593 1661 606
rect 1666 583 1669 606
rect 1234 533 1253 536
rect 1266 533 1277 536
rect 1290 533 1301 536
rect 1306 536 1309 546
rect 1314 543 1333 546
rect 1314 536 1317 543
rect 1306 533 1317 536
rect 1226 513 1229 526
rect 1234 503 1237 533
rect 1242 503 1245 516
rect 1218 413 1221 456
rect 1226 403 1229 446
rect 1234 413 1237 426
rect 1250 403 1253 516
rect 1258 413 1261 526
rect 1266 403 1269 526
rect 1274 443 1277 533
rect 1290 513 1293 526
rect 1298 493 1301 526
rect 1314 506 1317 533
rect 1322 523 1325 536
rect 1330 533 1333 543
rect 1338 523 1341 566
rect 1354 523 1357 546
rect 1362 523 1365 556
rect 1378 533 1381 546
rect 1314 503 1325 506
rect 1282 413 1285 436
rect 1290 403 1293 456
rect 1202 303 1205 336
rect 1210 333 1213 346
rect 1234 293 1237 326
rect 1258 323 1261 336
rect 1266 333 1269 356
rect 1306 353 1309 486
rect 1322 436 1325 503
rect 1386 456 1389 546
rect 1410 543 1413 556
rect 1394 506 1397 526
rect 1394 503 1401 506
rect 1378 453 1389 456
rect 1314 433 1325 436
rect 1314 413 1317 433
rect 1346 333 1349 386
rect 1354 346 1357 436
rect 1362 433 1373 436
rect 1362 413 1365 426
rect 1370 413 1373 433
rect 1354 343 1365 346
rect 1290 313 1293 326
rect 1322 313 1325 326
rect 1362 316 1365 343
rect 1370 323 1373 406
rect 1378 363 1381 453
rect 1398 426 1401 503
rect 1394 423 1401 426
rect 1386 403 1389 416
rect 1394 403 1397 423
rect 1410 406 1413 526
rect 1426 476 1429 536
rect 1434 533 1437 546
rect 1458 533 1469 536
rect 1418 473 1429 476
rect 1418 423 1421 473
rect 1434 446 1437 526
rect 1442 513 1445 526
rect 1434 443 1445 446
rect 1442 416 1445 443
rect 1450 423 1453 436
rect 1458 433 1461 533
rect 1466 513 1469 526
rect 1474 523 1477 546
rect 1482 533 1485 556
rect 1522 533 1533 536
rect 1554 533 1565 536
rect 1578 533 1581 546
rect 1522 526 1525 533
rect 1474 423 1477 436
rect 1410 403 1421 406
rect 1410 323 1413 336
rect 1362 313 1373 316
rect 1250 286 1253 306
rect 1386 293 1389 306
rect 1394 303 1397 316
rect 1418 313 1421 403
rect 1434 393 1437 416
rect 1442 413 1485 416
rect 1442 403 1445 413
rect 1482 403 1485 413
rect 1490 396 1493 526
rect 1498 513 1501 526
rect 1514 523 1525 526
rect 1506 413 1509 506
rect 1514 483 1517 516
rect 1522 433 1525 523
rect 1530 503 1533 526
rect 1562 513 1565 526
rect 1482 393 1493 396
rect 1498 393 1501 406
rect 1554 403 1557 426
rect 1482 366 1485 393
rect 1426 343 1429 366
rect 1482 363 1493 366
rect 1490 333 1493 363
rect 1562 326 1565 416
rect 1570 403 1573 506
rect 1578 476 1581 526
rect 1586 523 1589 536
rect 1594 503 1597 536
rect 1578 473 1589 476
rect 1586 423 1589 473
rect 1426 293 1429 326
rect 1546 323 1565 326
rect 1570 316 1573 396
rect 1578 323 1581 416
rect 1594 406 1597 486
rect 1618 436 1621 536
rect 1626 513 1629 526
rect 1634 493 1637 526
rect 1658 516 1661 546
rect 1650 513 1661 516
rect 1650 456 1653 513
rect 1650 453 1661 456
rect 1602 423 1605 436
rect 1610 433 1621 436
rect 1602 413 1613 416
rect 1594 403 1605 406
rect 1594 333 1597 366
rect 1602 343 1605 403
rect 1618 356 1621 426
rect 1610 353 1621 356
rect 1602 323 1605 336
rect 1562 313 1573 316
rect 1610 313 1613 353
rect 1618 333 1629 336
rect 1466 293 1469 306
rect 1250 283 1261 286
rect 1130 186 1133 206
rect 1138 193 1141 206
rect 1194 203 1197 216
rect 1218 213 1221 226
rect 1242 203 1245 276
rect 1258 226 1261 283
rect 1250 223 1261 226
rect 1250 203 1253 223
rect 1290 213 1293 256
rect 1322 213 1325 226
rect 1330 203 1333 266
rect 1378 233 1381 246
rect 1130 183 1149 186
rect 1058 113 1061 126
rect 1090 73 1093 136
rect 1138 133 1141 146
rect 1146 133 1149 183
rect 1114 103 1117 126
rect 1170 93 1173 126
rect 1194 103 1197 136
rect 1202 93 1205 166
rect 1250 133 1253 166
rect 1250 116 1253 126
rect 1258 123 1261 146
rect 1266 116 1269 196
rect 1274 133 1277 176
rect 1290 133 1293 146
rect 1298 123 1317 126
rect 1322 123 1325 136
rect 1250 113 1269 116
rect 1306 93 1309 116
rect 1314 103 1317 123
rect 1330 113 1333 126
rect 1338 103 1341 116
rect 1346 113 1349 166
rect 1354 113 1357 226
rect 1410 223 1421 226
rect 1442 223 1445 256
rect 1450 233 1477 236
rect 1410 213 1437 216
rect 1362 136 1365 146
rect 1362 133 1373 136
rect 1378 133 1381 196
rect 1402 146 1405 206
rect 1394 143 1405 146
rect 1386 123 1389 136
rect 1394 113 1397 143
rect 1418 133 1421 213
rect 1450 146 1453 226
rect 1474 206 1477 233
rect 1482 213 1485 236
rect 1490 213 1493 226
rect 1458 173 1461 206
rect 1474 203 1485 206
rect 1426 133 1429 146
rect 1434 143 1453 146
rect 1458 133 1461 166
rect 1498 156 1501 236
rect 1506 186 1509 256
rect 1522 223 1533 226
rect 1522 193 1525 216
rect 1530 213 1533 223
rect 1530 186 1533 206
rect 1562 203 1565 226
rect 1570 213 1573 236
rect 1586 213 1589 256
rect 1594 213 1597 226
rect 1586 193 1589 206
rect 1594 203 1605 206
rect 1506 183 1533 186
rect 1602 183 1605 203
rect 1482 153 1501 156
rect 1434 123 1445 126
rect 1466 123 1469 146
rect 1482 133 1485 153
rect 1618 146 1621 226
rect 1626 213 1629 256
rect 1626 183 1629 206
rect 1642 193 1645 416
rect 1650 333 1653 436
rect 1658 413 1661 453
rect 1666 373 1669 546
rect 1674 496 1677 666
rect 1682 593 1685 673
rect 1722 663 1725 683
rect 1690 616 1693 656
rect 1706 623 1725 626
rect 1690 613 1701 616
rect 1690 583 1693 606
rect 1698 593 1701 613
rect 1706 553 1709 623
rect 1722 613 1725 623
rect 1738 616 1741 786
rect 1738 613 1749 616
rect 1770 613 1773 806
rect 1778 803 1781 826
rect 1794 816 1797 966
rect 1818 853 1821 936
rect 1830 926 1833 973
rect 1842 933 1845 986
rect 1850 973 1853 1013
rect 1874 996 1877 1006
rect 1882 1003 1885 1056
rect 1890 996 1893 1016
rect 1874 993 1893 996
rect 1830 923 1837 926
rect 1778 706 1781 736
rect 1786 723 1789 816
rect 1794 813 1805 816
rect 1810 813 1813 826
rect 1778 703 1785 706
rect 1782 636 1785 703
rect 1778 633 1785 636
rect 1714 593 1717 606
rect 1722 583 1725 606
rect 1762 556 1765 576
rect 1754 553 1765 556
rect 1682 513 1685 526
rect 1674 493 1681 496
rect 1678 426 1681 493
rect 1690 466 1693 536
rect 1698 533 1701 546
rect 1714 483 1717 526
rect 1754 506 1757 553
rect 1770 513 1773 606
rect 1778 543 1781 633
rect 1786 573 1789 616
rect 1786 533 1789 566
rect 1794 533 1797 806
rect 1802 796 1805 806
rect 1818 803 1821 836
rect 1826 813 1829 866
rect 1826 796 1829 806
rect 1802 793 1829 796
rect 1818 733 1821 746
rect 1834 733 1837 923
rect 1842 793 1845 806
rect 1850 786 1853 816
rect 1858 803 1861 836
rect 1866 813 1869 926
rect 1890 896 1893 976
rect 1886 893 1893 896
rect 1866 793 1869 806
rect 1842 783 1853 786
rect 1842 733 1845 783
rect 1826 573 1829 646
rect 1834 613 1837 726
rect 1842 643 1845 726
rect 1850 723 1853 766
rect 1858 603 1861 746
rect 1866 723 1869 786
rect 1874 763 1877 846
rect 1886 806 1889 893
rect 1898 813 1901 1036
rect 1906 933 1909 1166
rect 1914 1083 1917 1146
rect 1914 916 1917 1016
rect 1910 913 1917 916
rect 1910 826 1913 913
rect 1910 823 1917 826
rect 1886 803 1893 806
rect 1842 533 1845 596
rect 1850 533 1853 576
rect 1874 553 1877 626
rect 1890 613 1893 803
rect 1914 793 1917 823
rect 1922 763 1925 1106
rect 1930 1003 1933 1096
rect 1930 893 1933 936
rect 1938 906 1941 1126
rect 1962 1113 1965 1186
rect 1970 1133 1973 1156
rect 1986 1153 1989 1236
rect 1994 1183 1997 1216
rect 2002 1153 2005 1526
rect 2050 1513 2053 1553
rect 2018 1466 2021 1486
rect 2014 1463 2021 1466
rect 2014 1376 2017 1463
rect 2014 1373 2021 1376
rect 2026 1373 2029 1476
rect 2034 1396 2037 1416
rect 2042 1403 2045 1416
rect 2050 1413 2053 1466
rect 2050 1396 2053 1406
rect 2034 1393 2053 1396
rect 2058 1386 2061 1583
rect 2066 1513 2069 1546
rect 2074 1483 2077 1566
rect 2082 1503 2085 1536
rect 2090 1533 2093 1646
rect 2098 1563 2101 1676
rect 2106 1603 2109 1626
rect 2114 1603 2117 1706
rect 2122 1703 2141 1706
rect 2162 1703 2165 1726
rect 2170 1696 2173 1806
rect 2178 1783 2181 1813
rect 2186 1713 2189 1806
rect 2194 1803 2197 1816
rect 2202 1796 2205 1866
rect 2210 1803 2213 1856
rect 2258 1836 2261 1936
rect 2274 1913 2277 1926
rect 2282 1896 2285 2006
rect 2290 1933 2293 2016
rect 2298 2013 2301 2123
rect 2314 2116 2317 2206
rect 2322 2126 2325 2243
rect 2354 2236 2357 2333
rect 2362 2313 2365 2326
rect 2450 2323 2453 2396
rect 2458 2383 2461 2396
rect 2466 2333 2469 2406
rect 2474 2403 2485 2406
rect 2474 2363 2477 2396
rect 2482 2373 2485 2403
rect 2498 2333 2501 2406
rect 2506 2326 2509 2506
rect 2514 2413 2517 2526
rect 2522 2383 2525 2536
rect 2530 2523 2533 2546
rect 2538 2533 2549 2536
rect 2538 2513 2541 2526
rect 2530 2423 2533 2456
rect 2546 2433 2549 2533
rect 2562 2513 2565 2526
rect 2362 2293 2365 2306
rect 2346 2233 2357 2236
rect 2346 2203 2349 2233
rect 2354 2213 2357 2226
rect 2362 2213 2365 2246
rect 2378 2243 2397 2246
rect 2378 2223 2381 2243
rect 2370 2213 2381 2216
rect 2386 2215 2389 2236
rect 2394 2206 2397 2243
rect 2410 2213 2413 2316
rect 2466 2313 2469 2326
rect 2498 2323 2509 2326
rect 2498 2313 2501 2323
rect 2418 2293 2421 2306
rect 2426 2303 2437 2306
rect 2450 2223 2453 2296
rect 2506 2256 2509 2316
rect 2514 2303 2517 2316
rect 2522 2303 2525 2326
rect 2530 2313 2533 2416
rect 2546 2413 2549 2426
rect 2562 2396 2565 2426
rect 2570 2403 2573 2426
rect 2594 2416 2597 2436
rect 2602 2423 2605 2436
rect 2578 2413 2589 2416
rect 2594 2413 2613 2416
rect 2554 2393 2565 2396
rect 2618 2396 2621 2406
rect 2626 2403 2629 2536
rect 2658 2416 2661 2436
rect 2618 2393 2629 2396
rect 2538 2333 2541 2386
rect 2554 2303 2557 2393
rect 2562 2303 2565 2376
rect 2506 2253 2517 2256
rect 2458 2223 2461 2236
rect 2474 2223 2477 2236
rect 2490 2233 2501 2236
rect 2490 2213 2493 2233
rect 2498 2213 2501 2226
rect 2506 2223 2509 2246
rect 2386 2203 2397 2206
rect 2330 2136 2333 2156
rect 2338 2143 2341 2196
rect 2386 2146 2389 2203
rect 2370 2143 2389 2146
rect 2394 2193 2413 2196
rect 2330 2133 2341 2136
rect 2322 2123 2333 2126
rect 2306 2113 2317 2116
rect 2306 2003 2309 2113
rect 2314 1933 2317 2106
rect 2322 2103 2325 2116
rect 2338 2106 2341 2133
rect 2334 2103 2341 2106
rect 2334 2026 2337 2103
rect 2322 2013 2325 2026
rect 2334 2023 2341 2026
rect 2338 2003 2341 2023
rect 2346 2013 2349 2126
rect 2354 2123 2357 2136
rect 2322 1923 2325 1996
rect 2354 1983 2357 2006
rect 2274 1893 2285 1896
rect 2258 1833 2269 1836
rect 2226 1813 2229 1826
rect 2258 1813 2261 1826
rect 2194 1793 2205 1796
rect 2162 1693 2173 1696
rect 2138 1613 2141 1626
rect 2066 1413 2069 1426
rect 2106 1413 2109 1426
rect 2018 1353 2021 1373
rect 2010 1323 2013 1336
rect 2018 1286 2021 1336
rect 2026 1313 2029 1326
rect 2018 1283 2029 1286
rect 2018 1206 2021 1276
rect 2026 1213 2029 1283
rect 2034 1256 2037 1386
rect 2050 1383 2061 1386
rect 2042 1303 2045 1356
rect 2034 1253 2045 1256
rect 2042 1213 2045 1253
rect 2010 1173 2013 1206
rect 2018 1203 2029 1206
rect 2018 1133 2021 1186
rect 2050 1183 2053 1383
rect 2066 1313 2069 1326
rect 2058 1203 2061 1216
rect 2026 1133 2029 1166
rect 2066 1153 2069 1306
rect 2074 1233 2077 1356
rect 2082 1313 2085 1406
rect 2114 1353 2117 1526
rect 2122 1363 2125 1516
rect 2114 1333 2117 1346
rect 2130 1333 2133 1496
rect 2138 1456 2141 1556
rect 2146 1513 2149 1536
rect 2138 1453 2149 1456
rect 2146 1383 2149 1453
rect 2154 1353 2157 1586
rect 2162 1493 2165 1693
rect 2170 1516 2173 1626
rect 2178 1533 2181 1606
rect 2194 1583 2197 1793
rect 2258 1783 2261 1806
rect 2218 1733 2229 1736
rect 2250 1733 2253 1746
rect 2266 1743 2269 1833
rect 2274 1803 2277 1893
rect 2290 1806 2293 1816
rect 2282 1803 2293 1806
rect 2282 1796 2285 1803
rect 2274 1793 2285 1796
rect 2202 1703 2205 1726
rect 2210 1693 2213 1706
rect 2218 1636 2221 1716
rect 2234 1713 2237 1726
rect 2242 1693 2245 1726
rect 2258 1703 2261 1716
rect 2266 1713 2269 1726
rect 2274 1703 2277 1793
rect 2290 1743 2293 1796
rect 2298 1793 2301 1806
rect 2330 1763 2333 1816
rect 2338 1813 2341 1826
rect 2346 1803 2349 1946
rect 2362 1876 2365 2036
rect 2370 2013 2373 2143
rect 2378 2123 2381 2136
rect 2386 2123 2389 2136
rect 2394 2133 2397 2193
rect 2378 2103 2381 2116
rect 2402 2103 2405 2146
rect 2410 2143 2413 2156
rect 2482 2153 2485 2206
rect 2514 2176 2517 2253
rect 2522 2216 2525 2226
rect 2522 2213 2533 2216
rect 2562 2213 2565 2226
rect 2578 2213 2581 2316
rect 2586 2246 2589 2336
rect 2650 2333 2653 2416
rect 2658 2413 2665 2416
rect 2662 2346 2665 2413
rect 2658 2343 2665 2346
rect 2658 2316 2661 2343
rect 2650 2313 2661 2316
rect 2650 2246 2653 2313
rect 2586 2243 2605 2246
rect 2650 2243 2661 2246
rect 2490 2173 2517 2176
rect 2530 2176 2533 2213
rect 2586 2203 2589 2236
rect 2554 2183 2565 2186
rect 2530 2173 2549 2176
rect 2410 2123 2413 2136
rect 2490 2133 2493 2173
rect 2514 2163 2517 2173
rect 2498 2133 2501 2146
rect 2546 2133 2549 2173
rect 2378 2006 2381 2026
rect 2370 2003 2381 2006
rect 2386 1943 2389 2006
rect 2426 1936 2429 1946
rect 2386 1933 2397 1936
rect 2402 1933 2429 1936
rect 2378 1923 2397 1926
rect 2362 1873 2373 1876
rect 2354 1803 2365 1806
rect 2370 1803 2373 1873
rect 2386 1813 2389 1916
rect 2402 1903 2405 1916
rect 2410 1913 2421 1916
rect 2402 1813 2405 1826
rect 2418 1813 2421 1836
rect 2426 1803 2429 1816
rect 2346 1746 2349 1776
rect 2354 1753 2357 1803
rect 2362 1773 2365 1796
rect 2346 1743 2357 1746
rect 2290 1723 2293 1736
rect 2202 1633 2221 1636
rect 2202 1603 2205 1633
rect 2226 1613 2229 1626
rect 2258 1566 2261 1626
rect 2266 1583 2269 1616
rect 2274 1603 2277 1616
rect 2282 1613 2285 1716
rect 2314 1623 2317 1726
rect 2322 1683 2325 1726
rect 2338 1716 2341 1736
rect 2354 1733 2357 1743
rect 2354 1716 2357 1726
rect 2338 1713 2357 1716
rect 2282 1573 2285 1606
rect 2234 1536 2237 1566
rect 2258 1563 2301 1566
rect 2226 1533 2237 1536
rect 2242 1533 2245 1546
rect 2250 1533 2253 1556
rect 2170 1513 2177 1516
rect 2202 1513 2205 1526
rect 2226 1513 2229 1526
rect 2174 1446 2177 1513
rect 2234 1476 2237 1533
rect 2162 1413 2165 1446
rect 2170 1443 2177 1446
rect 2226 1473 2237 1476
rect 2170 1413 2173 1443
rect 2194 1413 2197 1436
rect 2162 1403 2173 1406
rect 2218 1403 2221 1416
rect 2226 1403 2229 1473
rect 2258 1413 2261 1466
rect 2274 1403 2277 1456
rect 2282 1403 2285 1446
rect 2298 1413 2301 1563
rect 2306 1533 2309 1586
rect 2330 1563 2333 1616
rect 2338 1603 2341 1706
rect 2362 1703 2365 1766
rect 2378 1733 2381 1746
rect 2386 1743 2389 1776
rect 2386 1726 2389 1736
rect 2370 1723 2389 1726
rect 2354 1633 2357 1686
rect 2346 1606 2349 1626
rect 2362 1613 2365 1636
rect 2370 1623 2373 1723
rect 2394 1633 2397 1756
rect 2426 1733 2429 1786
rect 2434 1773 2437 2046
rect 2442 2023 2445 2036
rect 2466 2023 2469 2126
rect 2474 2023 2493 2026
rect 2442 2013 2469 2016
rect 2458 1946 2461 2006
rect 2466 2003 2469 2013
rect 2458 1943 2469 1946
rect 2474 1936 2477 2023
rect 2490 1946 2493 2006
rect 2498 2003 2501 2126
rect 2530 2013 2533 2026
rect 2546 2013 2549 2126
rect 2426 1703 2429 1716
rect 2434 1636 2437 1756
rect 2442 1723 2445 1816
rect 2450 1813 2453 1936
rect 2458 1933 2477 1936
rect 2482 1943 2493 1946
rect 2458 1903 2461 1933
rect 2466 1913 2469 1926
rect 2482 1916 2485 1943
rect 2498 1926 2501 1996
rect 2474 1913 2485 1916
rect 2494 1923 2501 1926
rect 2474 1896 2477 1913
rect 2470 1893 2477 1896
rect 2470 1826 2473 1893
rect 2470 1823 2477 1826
rect 2482 1823 2485 1906
rect 2494 1856 2497 1923
rect 2506 1866 2509 1946
rect 2530 1933 2533 1986
rect 2546 1946 2549 2006
rect 2554 1976 2557 2183
rect 2594 2153 2597 2216
rect 2602 2133 2605 2243
rect 2602 2113 2605 2126
rect 2610 2106 2613 2166
rect 2658 2146 2661 2243
rect 2666 2153 2669 2326
rect 2658 2143 2669 2146
rect 2602 2103 2613 2106
rect 2578 2013 2581 2046
rect 2602 2013 2605 2103
rect 2554 1973 2573 1976
rect 2546 1943 2557 1946
rect 2506 1863 2513 1866
rect 2494 1853 2501 1856
rect 2458 1803 2469 1806
rect 2474 1793 2477 1823
rect 2450 1733 2477 1736
rect 2378 1613 2381 1626
rect 2394 1613 2397 1626
rect 2402 1613 2405 1636
rect 2434 1633 2445 1636
rect 2450 1633 2453 1726
rect 2346 1603 2357 1606
rect 2354 1533 2357 1603
rect 2322 1486 2325 1526
rect 2330 1496 2333 1526
rect 2354 1503 2357 1526
rect 2330 1493 2345 1496
rect 2322 1483 2333 1486
rect 2306 1413 2309 1426
rect 2330 1403 2333 1483
rect 2242 1383 2253 1386
rect 2090 1213 2093 1226
rect 1986 1033 1989 1126
rect 1946 1013 1949 1026
rect 1970 1013 1973 1026
rect 1994 933 1997 1126
rect 2018 1113 2021 1126
rect 2002 973 2005 1036
rect 2010 933 2013 1106
rect 2074 1063 2077 1136
rect 2082 1133 2085 1166
rect 2114 1163 2117 1326
rect 2122 1153 2125 1226
rect 2130 1133 2133 1326
rect 2146 1273 2149 1326
rect 2178 1303 2181 1336
rect 2138 1213 2141 1246
rect 2138 1183 2141 1206
rect 2138 1133 2141 1166
rect 2018 1003 2021 1046
rect 2034 953 2037 1036
rect 2082 1033 2085 1126
rect 2098 1073 2101 1126
rect 2106 1033 2109 1126
rect 2146 1106 2149 1216
rect 2154 1213 2157 1226
rect 2154 1203 2165 1206
rect 2154 1123 2157 1146
rect 2162 1133 2165 1203
rect 2170 1133 2173 1146
rect 2178 1126 2181 1276
rect 2186 1223 2189 1336
rect 2194 1313 2197 1326
rect 2210 1306 2213 1336
rect 2234 1313 2237 1326
rect 2202 1303 2213 1306
rect 2202 1276 2205 1303
rect 2202 1273 2213 1276
rect 2210 1216 2213 1273
rect 2202 1213 2213 1216
rect 2170 1123 2181 1126
rect 2122 1103 2149 1106
rect 2058 1013 2061 1026
rect 2090 1013 2093 1026
rect 2042 966 2045 1006
rect 2042 963 2061 966
rect 2058 933 2061 963
rect 2066 933 2069 946
rect 1938 903 1949 906
rect 1930 776 1933 816
rect 1938 803 1941 816
rect 1946 813 1949 903
rect 1954 806 1957 876
rect 1962 863 1965 926
rect 1946 793 1949 806
rect 1954 803 1965 806
rect 1930 773 1949 776
rect 1930 733 1933 746
rect 1946 733 1949 773
rect 1906 713 1909 726
rect 1946 713 1949 726
rect 1898 613 1901 626
rect 1922 576 1925 626
rect 1930 593 1933 616
rect 1962 613 1965 803
rect 1994 796 1997 816
rect 2002 803 2005 816
rect 2018 813 2021 826
rect 2010 796 2013 806
rect 1994 793 2013 796
rect 2026 786 2029 816
rect 2018 783 2029 786
rect 2034 783 2037 806
rect 2042 786 2045 926
rect 2074 923 2077 956
rect 2066 813 2069 826
rect 2090 813 2093 1006
rect 2098 1003 2101 1016
rect 2106 963 2109 1006
rect 2114 953 2117 1016
rect 2122 933 2125 1103
rect 2130 1013 2133 1046
rect 2130 953 2133 1006
rect 2138 1003 2141 1056
rect 2146 1013 2149 1026
rect 2154 933 2157 966
rect 2042 783 2069 786
rect 1994 703 1997 766
rect 2018 723 2021 783
rect 2042 723 2045 746
rect 2058 723 2061 776
rect 2066 696 2069 783
rect 2090 706 2093 806
rect 2098 773 2101 816
rect 2106 813 2109 886
rect 2106 723 2109 756
rect 2114 723 2117 816
rect 2122 813 2125 926
rect 2130 906 2133 926
rect 2130 903 2137 906
rect 2134 836 2137 903
rect 2146 883 2149 926
rect 2162 836 2165 1076
rect 2170 1053 2173 1123
rect 2186 1113 2189 1126
rect 2202 1073 2205 1213
rect 2226 1113 2229 1126
rect 2186 1013 2189 1026
rect 2170 903 2173 966
rect 2202 956 2205 1026
rect 2178 953 2205 956
rect 2226 953 2229 1036
rect 2130 833 2137 836
rect 2146 833 2165 836
rect 2130 813 2133 833
rect 2130 783 2133 806
rect 2138 743 2141 816
rect 2146 753 2149 833
rect 2138 723 2141 736
rect 2090 703 2101 706
rect 2058 693 2069 696
rect 1906 573 1925 576
rect 1898 533 1901 556
rect 1906 533 1909 573
rect 1938 563 1941 606
rect 1754 503 1765 506
rect 1690 463 1701 466
rect 1674 423 1681 426
rect 1674 403 1677 423
rect 1698 396 1701 463
rect 1690 393 1701 396
rect 1658 343 1685 346
rect 1666 333 1677 336
rect 1682 333 1685 343
rect 1690 336 1693 393
rect 1690 333 1701 336
rect 1650 313 1653 326
rect 1658 293 1661 326
rect 1682 306 1685 326
rect 1690 313 1693 326
rect 1698 306 1701 333
rect 1706 313 1709 326
rect 1714 323 1717 336
rect 1722 333 1725 496
rect 1762 423 1765 503
rect 1778 413 1781 426
rect 1786 413 1789 436
rect 1810 413 1813 526
rect 1778 403 1789 406
rect 1770 333 1773 376
rect 1746 323 1757 326
rect 1682 303 1701 306
rect 1770 263 1773 326
rect 1778 316 1781 396
rect 1834 393 1837 406
rect 1842 383 1845 426
rect 1810 333 1813 376
rect 1850 356 1853 526
rect 1842 353 1853 356
rect 1778 313 1797 316
rect 1650 223 1653 236
rect 1490 143 1501 146
rect 1610 143 1621 146
rect 1498 133 1509 136
rect 1362 103 1373 106
rect 1490 103 1493 126
rect 1514 123 1517 136
rect 1610 133 1613 143
rect 1618 133 1629 136
rect 1546 103 1549 126
rect 1578 103 1581 126
rect 1634 103 1637 126
rect 1650 123 1653 216
rect 1658 146 1661 226
rect 1666 223 1669 236
rect 1674 193 1677 216
rect 1682 213 1685 226
rect 1698 203 1701 216
rect 1658 143 1677 146
rect 1674 113 1677 143
rect 1682 133 1685 146
rect 1682 103 1685 116
rect 1706 113 1709 216
rect 1714 213 1717 246
rect 1730 203 1733 216
rect 1714 193 1733 196
rect 1722 133 1725 186
rect 1730 133 1733 193
rect 1746 183 1749 236
rect 1794 226 1797 313
rect 1778 223 1797 226
rect 1770 186 1773 196
rect 1778 193 1781 223
rect 1818 203 1821 346
rect 1826 313 1829 346
rect 1842 296 1845 353
rect 1850 326 1853 346
rect 1858 336 1861 436
rect 1866 343 1869 436
rect 1874 383 1877 526
rect 1898 513 1901 526
rect 1954 506 1957 526
rect 1882 376 1885 416
rect 1874 373 1885 376
rect 1874 363 1877 373
rect 1890 363 1893 406
rect 1898 403 1901 506
rect 1946 503 1957 506
rect 1986 503 1989 616
rect 2018 613 2021 626
rect 1994 593 1997 606
rect 2058 566 2061 693
rect 2058 563 2069 566
rect 2010 533 2013 546
rect 2018 513 2021 556
rect 1946 403 1949 503
rect 1858 333 1869 336
rect 1850 323 1861 326
rect 1858 313 1861 323
rect 1834 293 1845 296
rect 1834 236 1837 293
rect 1834 233 1845 236
rect 1842 213 1845 233
rect 1850 213 1853 306
rect 1866 213 1869 333
rect 1890 313 1893 326
rect 1898 306 1901 386
rect 1946 343 1949 366
rect 1890 303 1901 306
rect 1890 233 1893 303
rect 1906 256 1909 326
rect 1922 303 1925 326
rect 1930 323 1933 336
rect 1954 333 1957 426
rect 1962 413 1965 436
rect 1970 416 1973 436
rect 1978 423 1981 466
rect 2050 436 2053 506
rect 1970 413 1989 416
rect 2002 406 2005 416
rect 2018 413 2021 436
rect 2034 433 2053 436
rect 1978 403 2005 406
rect 1962 333 1965 366
rect 1898 253 1909 256
rect 1834 203 1853 206
rect 1826 193 1845 196
rect 1850 193 1853 203
rect 1770 183 1781 186
rect 1722 113 1725 126
rect 1730 123 1749 126
rect 1762 123 1765 136
rect 1770 123 1773 136
rect 1778 133 1781 183
rect 1842 133 1845 193
rect 1818 123 1829 126
rect 1890 123 1893 216
rect 1898 133 1901 253
rect 1954 236 1957 326
rect 1970 323 1973 346
rect 1978 336 1981 403
rect 1986 346 1989 396
rect 2034 363 2037 433
rect 1986 343 1997 346
rect 2026 343 2029 356
rect 1978 333 1989 336
rect 1994 326 1997 343
rect 2042 336 2045 426
rect 2058 383 2061 436
rect 2066 396 2069 563
rect 2074 403 2077 546
rect 2082 433 2085 686
rect 2098 616 2101 703
rect 2146 676 2149 706
rect 2138 673 2149 676
rect 2122 623 2125 636
rect 2094 613 2101 616
rect 2138 616 2141 673
rect 2154 623 2157 816
rect 2162 733 2165 826
rect 2138 613 2149 616
rect 2094 556 2097 613
rect 2090 553 2097 556
rect 2090 503 2093 553
rect 2098 523 2101 536
rect 2106 533 2109 596
rect 2098 413 2101 516
rect 2114 506 2117 526
rect 2122 513 2125 546
rect 2138 513 2141 526
rect 2114 503 2133 506
rect 2106 413 2109 426
rect 2122 403 2125 426
rect 2066 393 2077 396
rect 2130 393 2133 436
rect 2146 413 2149 613
rect 2162 603 2165 726
rect 2170 613 2173 746
rect 2178 683 2181 953
rect 2234 933 2237 1216
rect 2242 1013 2245 1376
rect 2250 1366 2253 1383
rect 2274 1376 2277 1396
rect 2274 1373 2281 1376
rect 2250 1363 2257 1366
rect 2254 1176 2257 1363
rect 2278 1286 2281 1373
rect 2274 1283 2281 1286
rect 2274 1236 2277 1283
rect 2290 1243 2293 1386
rect 2342 1366 2345 1493
rect 2298 1333 2301 1366
rect 2342 1363 2349 1366
rect 2298 1236 2301 1326
rect 2346 1306 2349 1363
rect 2250 1173 2257 1176
rect 2266 1233 2277 1236
rect 2282 1233 2301 1236
rect 2330 1303 2349 1306
rect 2250 986 2253 1173
rect 2266 1123 2269 1233
rect 2274 1203 2277 1216
rect 2282 1213 2285 1233
rect 2330 1183 2333 1303
rect 2354 1223 2357 1466
rect 2274 1093 2277 1146
rect 2282 1123 2285 1166
rect 2338 1133 2341 1206
rect 2346 1193 2349 1216
rect 2362 1213 2365 1576
rect 2370 1496 2373 1606
rect 2434 1573 2437 1626
rect 2378 1513 2381 1546
rect 2386 1523 2389 1536
rect 2442 1533 2445 1633
rect 2458 1616 2461 1716
rect 2474 1713 2477 1733
rect 2482 1723 2485 1816
rect 2490 1753 2493 1836
rect 2498 1783 2501 1853
rect 2510 1776 2513 1863
rect 2498 1746 2501 1776
rect 2490 1743 2501 1746
rect 2506 1773 2513 1776
rect 2506 1743 2509 1773
rect 2522 1756 2525 1916
rect 2530 1813 2533 1836
rect 2538 1813 2541 1936
rect 2554 1866 2557 1943
rect 2546 1863 2557 1866
rect 2546 1833 2549 1863
rect 2570 1846 2573 1973
rect 2602 1926 2605 2006
rect 2610 1976 2613 2016
rect 2634 2013 2637 2126
rect 2642 2013 2645 2026
rect 2658 2013 2661 2136
rect 2666 2113 2669 2143
rect 2658 1976 2661 2006
rect 2610 1973 2629 1976
rect 2602 1923 2613 1926
rect 2554 1843 2573 1846
rect 2546 1803 2549 1826
rect 2514 1753 2541 1756
rect 2466 1693 2469 1706
rect 2482 1683 2485 1716
rect 2490 1666 2493 1736
rect 2486 1663 2493 1666
rect 2466 1623 2469 1636
rect 2450 1613 2461 1616
rect 2474 1613 2477 1626
rect 2486 1576 2489 1663
rect 2498 1613 2501 1736
rect 2498 1596 2501 1606
rect 2506 1603 2509 1726
rect 2514 1683 2517 1753
rect 2522 1716 2525 1746
rect 2530 1723 2533 1736
rect 2538 1733 2541 1753
rect 2538 1716 2541 1726
rect 2522 1713 2541 1716
rect 2514 1596 2517 1646
rect 2546 1643 2549 1736
rect 2554 1716 2557 1843
rect 2562 1733 2565 1806
rect 2570 1783 2573 1806
rect 2578 1746 2581 1816
rect 2586 1803 2589 1826
rect 2594 1813 2597 1916
rect 2610 1876 2613 1923
rect 2602 1873 2613 1876
rect 2602 1823 2605 1873
rect 2626 1856 2629 1973
rect 2610 1853 2629 1856
rect 2650 1973 2661 1976
rect 2570 1733 2573 1746
rect 2578 1743 2589 1746
rect 2586 1723 2589 1743
rect 2554 1713 2561 1716
rect 2558 1646 2561 1713
rect 2570 1703 2573 1716
rect 2594 1693 2597 1806
rect 2602 1803 2605 1816
rect 2602 1783 2605 1796
rect 2602 1703 2605 1716
rect 2554 1643 2561 1646
rect 2522 1613 2525 1636
rect 2498 1593 2525 1596
rect 2486 1573 2493 1576
rect 2370 1493 2381 1496
rect 2266 1013 2269 1026
rect 2298 1013 2301 1066
rect 2306 1006 2309 1126
rect 2314 1096 2317 1126
rect 2346 1116 2349 1156
rect 2338 1113 2349 1116
rect 2354 1113 2357 1206
rect 2370 1136 2373 1426
rect 2378 1343 2381 1493
rect 2386 1343 2389 1406
rect 2378 1203 2381 1336
rect 2386 1303 2389 1316
rect 2394 1243 2397 1436
rect 2402 1413 2405 1506
rect 2410 1476 2413 1526
rect 2418 1493 2421 1516
rect 2426 1513 2429 1526
rect 2434 1523 2461 1526
rect 2434 1513 2437 1523
rect 2410 1473 2421 1476
rect 2362 1133 2373 1136
rect 2338 1096 2341 1113
rect 2314 1093 2325 1096
rect 2298 1003 2309 1006
rect 2250 983 2261 986
rect 2242 946 2245 976
rect 2242 943 2253 946
rect 2258 943 2261 983
rect 2322 966 2325 1093
rect 2334 1093 2341 1096
rect 2334 1006 2337 1093
rect 2346 1013 2349 1106
rect 2362 1046 2365 1133
rect 2370 1113 2373 1126
rect 2370 1063 2373 1106
rect 2378 1103 2381 1116
rect 2386 1106 2389 1226
rect 2394 1123 2397 1236
rect 2402 1153 2405 1346
rect 2410 1303 2413 1316
rect 2418 1313 2421 1473
rect 2442 1413 2445 1516
rect 2450 1503 2453 1516
rect 2458 1513 2461 1523
rect 2466 1503 2469 1526
rect 2426 1306 2429 1346
rect 2434 1333 2437 1396
rect 2418 1303 2429 1306
rect 2402 1133 2405 1146
rect 2410 1116 2413 1246
rect 2402 1113 2413 1116
rect 2386 1103 2397 1106
rect 2386 1083 2389 1096
rect 2394 1076 2397 1103
rect 2378 1073 2397 1076
rect 2362 1043 2373 1046
rect 2354 1033 2365 1036
rect 2334 1003 2341 1006
rect 2314 963 2325 966
rect 2186 913 2189 926
rect 2210 913 2213 926
rect 2186 733 2189 756
rect 2194 703 2197 886
rect 2218 813 2221 826
rect 2202 633 2205 716
rect 2218 713 2221 756
rect 2210 693 2213 706
rect 2194 613 2197 626
rect 2226 623 2229 836
rect 2234 703 2237 826
rect 2242 823 2245 936
rect 2250 883 2253 943
rect 2250 816 2253 836
rect 2258 823 2261 926
rect 2242 813 2253 816
rect 2266 813 2269 936
rect 2274 833 2277 936
rect 2298 933 2301 946
rect 2274 813 2277 826
rect 2242 783 2245 806
rect 2282 796 2285 926
rect 2306 916 2309 956
rect 2302 913 2309 916
rect 2290 803 2293 846
rect 2302 826 2305 913
rect 2314 836 2317 963
rect 2338 953 2341 1003
rect 2354 993 2357 1026
rect 2362 1013 2365 1033
rect 2362 943 2365 1006
rect 2330 903 2333 926
rect 2362 913 2365 936
rect 2314 833 2325 836
rect 2298 823 2305 826
rect 2298 803 2301 823
rect 2282 793 2293 796
rect 2242 733 2269 736
rect 2274 733 2285 736
rect 2234 613 2237 646
rect 2242 613 2245 733
rect 2258 723 2269 726
rect 2178 513 2181 606
rect 2250 603 2253 616
rect 2258 596 2261 716
rect 2266 713 2269 723
rect 2282 643 2285 726
rect 2250 593 2261 596
rect 2178 403 2181 416
rect 2186 403 2189 526
rect 2250 513 2253 593
rect 2258 506 2261 566
rect 2266 513 2269 616
rect 2274 593 2277 636
rect 2274 543 2277 556
rect 2290 543 2293 793
rect 2306 746 2309 816
rect 2314 813 2317 826
rect 2322 746 2325 833
rect 2346 756 2349 816
rect 2354 803 2357 906
rect 2362 813 2365 826
rect 2346 753 2357 756
rect 2302 743 2309 746
rect 2314 743 2325 746
rect 2302 636 2305 743
rect 2314 693 2317 743
rect 2322 713 2325 736
rect 2298 633 2305 636
rect 2258 503 2269 506
rect 2210 413 2213 436
rect 2234 393 2237 406
rect 2242 403 2245 436
rect 2266 413 2269 503
rect 2290 496 2293 516
rect 2298 503 2301 633
rect 2290 493 2301 496
rect 2298 423 2301 493
rect 2290 403 2293 416
rect 2306 413 2309 616
rect 2322 603 2325 626
rect 2330 543 2333 726
rect 2338 723 2341 736
rect 2338 526 2341 716
rect 2346 713 2349 746
rect 2354 723 2357 753
rect 2362 723 2365 806
rect 2362 703 2365 716
rect 2370 696 2373 1043
rect 2378 1003 2381 1073
rect 2386 1003 2389 1016
rect 2394 996 2397 1066
rect 2378 943 2381 996
rect 2386 993 2397 996
rect 2386 936 2389 993
rect 2378 933 2389 936
rect 2386 906 2389 926
rect 2382 903 2389 906
rect 2382 836 2385 903
rect 2382 833 2389 836
rect 2378 733 2381 816
rect 2386 723 2389 833
rect 2394 803 2397 916
rect 2394 733 2397 776
rect 2402 713 2405 1113
rect 2418 1106 2421 1303
rect 2434 1226 2437 1256
rect 2442 1233 2445 1346
rect 2450 1253 2453 1396
rect 2458 1366 2461 1416
rect 2466 1403 2469 1496
rect 2474 1413 2477 1526
rect 2482 1503 2485 1556
rect 2482 1413 2485 1426
rect 2458 1363 2469 1366
rect 2458 1343 2461 1356
rect 2466 1336 2469 1363
rect 2466 1333 2477 1336
rect 2458 1303 2461 1326
rect 2466 1313 2469 1326
rect 2426 1213 2429 1226
rect 2434 1223 2445 1226
rect 2426 1163 2429 1206
rect 2434 1143 2437 1206
rect 2442 1203 2445 1223
rect 2450 1213 2453 1226
rect 2474 1213 2477 1333
rect 2482 1303 2485 1336
rect 2466 1203 2477 1206
rect 2482 1193 2485 1206
rect 2426 1113 2429 1126
rect 2434 1113 2437 1126
rect 2410 1103 2421 1106
rect 2410 1076 2413 1096
rect 2450 1083 2453 1166
rect 2458 1126 2461 1146
rect 2458 1123 2465 1126
rect 2462 1076 2465 1123
rect 2474 1093 2477 1146
rect 2482 1133 2485 1156
rect 2410 1073 2417 1076
rect 2414 956 2417 1073
rect 2458 1073 2465 1076
rect 2458 1026 2461 1073
rect 2474 1026 2477 1086
rect 2426 1023 2461 1026
rect 2466 1023 2477 1026
rect 2442 973 2445 1016
rect 2466 1006 2469 1023
rect 2450 1003 2469 1006
rect 2450 983 2453 1003
rect 2474 963 2477 1006
rect 2410 953 2417 956
rect 2410 903 2413 953
rect 2426 876 2429 956
rect 2434 923 2437 936
rect 2482 933 2485 1026
rect 2422 873 2429 876
rect 2422 826 2425 873
rect 2330 523 2341 526
rect 2314 433 2317 516
rect 2330 446 2333 523
rect 2346 456 2349 696
rect 2362 693 2373 696
rect 2354 553 2357 616
rect 2346 453 2353 456
rect 2330 443 2341 446
rect 2322 413 2325 426
rect 2330 403 2333 416
rect 2026 326 2029 336
rect 1938 233 1957 236
rect 1938 203 1941 233
rect 1922 123 1933 126
rect 1954 113 1957 226
rect 1970 213 1973 226
rect 1978 213 1981 326
rect 1986 323 1997 326
rect 2010 323 2029 326
rect 2034 333 2045 336
rect 2050 333 2053 376
rect 2034 323 2037 333
rect 1986 213 1989 323
rect 1994 313 2005 316
rect 2010 303 2013 323
rect 2018 313 2029 316
rect 2018 293 2021 306
rect 1994 223 1997 236
rect 2026 226 2029 313
rect 2042 246 2045 326
rect 2050 313 2053 326
rect 2042 243 2053 246
rect 2058 243 2061 356
rect 2066 313 2069 366
rect 1978 203 1989 206
rect 2002 133 2005 146
rect 2010 123 2013 216
rect 2018 213 2021 226
rect 2026 223 2037 226
rect 2042 223 2045 236
rect 2026 203 2029 216
rect 2034 156 2037 223
rect 2050 206 2053 243
rect 2050 203 2061 206
rect 2018 153 2037 156
rect 2018 133 2021 153
rect 2026 133 2029 146
rect 2034 133 2037 153
rect 2066 133 2069 236
rect 2074 223 2077 393
rect 2082 333 2085 386
rect 2082 313 2085 326
rect 2090 323 2093 336
rect 2098 303 2101 346
rect 2106 286 2109 336
rect 2114 313 2117 326
rect 2098 283 2109 286
rect 2074 193 2077 206
rect 2082 203 2093 206
rect 2090 183 2093 203
rect 2098 143 2101 283
rect 2122 256 2125 386
rect 2130 333 2133 346
rect 2138 273 2141 326
rect 2210 296 2213 346
rect 2218 303 2221 316
rect 2210 293 2221 296
rect 2114 253 2125 256
rect 2106 213 2109 246
rect 2114 206 2117 253
rect 2122 213 2125 226
rect 2106 203 2117 206
rect 2106 193 2109 203
rect 2122 183 2125 206
rect 2170 203 2173 246
rect 2178 153 2181 226
rect 2194 156 2197 236
rect 2202 233 2213 236
rect 2202 213 2205 226
rect 2210 213 2213 233
rect 2194 153 2205 156
rect 2106 133 2117 136
rect 2114 113 2125 116
rect 2202 113 2205 153
rect 2210 103 2213 206
rect 2218 183 2221 293
rect 2226 223 2229 236
rect 2242 233 2245 346
rect 2250 333 2285 336
rect 2250 313 2253 326
rect 2258 293 2261 326
rect 2266 236 2269 316
rect 2282 306 2285 333
rect 2290 313 2293 386
rect 2338 383 2341 443
rect 2350 386 2353 453
rect 2362 396 2365 693
rect 2410 603 2413 826
rect 2422 823 2429 826
rect 2434 823 2437 866
rect 2466 826 2469 906
rect 2466 823 2477 826
rect 2482 823 2485 926
rect 2426 803 2429 823
rect 2450 756 2453 816
rect 2466 803 2469 823
rect 2434 753 2453 756
rect 2418 733 2429 736
rect 2418 603 2421 626
rect 2370 533 2373 546
rect 2378 533 2381 556
rect 2370 506 2373 526
rect 2370 503 2381 506
rect 2378 446 2381 503
rect 2370 443 2381 446
rect 2370 403 2373 443
rect 2378 423 2389 426
rect 2362 393 2373 396
rect 2346 383 2353 386
rect 2306 333 2317 336
rect 2330 333 2333 346
rect 2250 223 2253 236
rect 2258 233 2269 236
rect 2274 303 2285 306
rect 2274 233 2277 303
rect 2226 213 2245 216
rect 2226 123 2229 213
rect 2258 193 2261 233
rect 2282 226 2285 296
rect 2290 283 2293 306
rect 2298 293 2301 326
rect 2314 313 2317 326
rect 2330 303 2333 326
rect 2338 323 2341 336
rect 2282 223 2293 226
rect 2266 186 2269 206
rect 2258 183 2269 186
rect 2258 146 2261 183
rect 2274 163 2277 206
rect 2282 203 2285 216
rect 2234 143 2261 146
rect 2234 133 2237 143
rect 2242 133 2253 136
rect 2258 116 2261 126
rect 2266 123 2277 126
rect 2258 113 2269 116
rect 2282 103 2285 176
rect 2290 133 2293 223
rect 2314 213 2325 216
rect 2330 213 2333 286
rect 2346 283 2349 383
rect 2370 356 2373 393
rect 2370 353 2381 356
rect 2370 333 2373 353
rect 2378 333 2381 346
rect 2386 343 2389 396
rect 2362 236 2365 326
rect 2386 306 2389 336
rect 2394 313 2397 586
rect 2426 583 2429 726
rect 2434 723 2437 753
rect 2442 716 2445 746
rect 2490 733 2493 1573
rect 2498 1333 2501 1546
rect 2514 1536 2517 1586
rect 2530 1553 2533 1606
rect 2538 1583 2541 1606
rect 2546 1603 2549 1616
rect 2546 1553 2549 1596
rect 2522 1543 2549 1546
rect 2506 1533 2517 1536
rect 2506 1483 2509 1533
rect 2514 1513 2517 1526
rect 2498 1313 2501 1326
rect 2506 1306 2509 1406
rect 2514 1403 2517 1426
rect 2522 1393 2525 1536
rect 2530 1413 2533 1426
rect 2538 1403 2541 1536
rect 2546 1533 2549 1543
rect 2554 1513 2557 1643
rect 2578 1613 2581 1686
rect 2586 1613 2589 1626
rect 2562 1523 2565 1586
rect 2514 1333 2517 1356
rect 2546 1336 2549 1486
rect 2562 1413 2565 1426
rect 2554 1403 2565 1406
rect 2570 1396 2573 1516
rect 2586 1413 2589 1526
rect 2594 1523 2597 1586
rect 2602 1573 2605 1686
rect 2610 1613 2613 1853
rect 2650 1846 2653 1973
rect 2650 1843 2661 1846
rect 2618 1826 2621 1836
rect 2618 1823 2637 1826
rect 2618 1813 2621 1823
rect 2618 1726 2621 1806
rect 2626 1783 2629 1816
rect 2634 1733 2637 1823
rect 2642 1806 2645 1826
rect 2642 1803 2649 1806
rect 2618 1723 2629 1726
rect 2626 1703 2629 1723
rect 2634 1613 2637 1716
rect 2646 1706 2649 1803
rect 2642 1703 2649 1706
rect 2642 1683 2645 1703
rect 2602 1533 2605 1566
rect 2610 1543 2613 1606
rect 2658 1596 2661 1843
rect 2666 1603 2669 2006
rect 2658 1593 2669 1596
rect 2594 1486 2597 1506
rect 2610 1503 2613 1536
rect 2594 1483 2605 1486
rect 2602 1426 2605 1483
rect 2594 1423 2605 1426
rect 2562 1393 2573 1396
rect 2546 1333 2557 1336
rect 2562 1326 2565 1393
rect 2594 1353 2597 1423
rect 2522 1323 2541 1326
rect 2498 1303 2509 1306
rect 2498 1223 2501 1303
rect 2514 1246 2517 1316
rect 2522 1303 2525 1316
rect 2506 1243 2517 1246
rect 2498 1146 2501 1206
rect 2506 1193 2509 1243
rect 2514 1233 2533 1236
rect 2514 1203 2517 1233
rect 2522 1223 2533 1226
rect 2522 1193 2525 1206
rect 2498 1143 2509 1146
rect 2498 1123 2501 1136
rect 2506 1123 2509 1143
rect 2514 1123 2517 1176
rect 2530 1163 2533 1223
rect 2538 1213 2541 1256
rect 2546 1233 2549 1326
rect 2554 1323 2565 1326
rect 2570 1323 2573 1336
rect 2554 1223 2557 1323
rect 2570 1303 2573 1316
rect 2578 1313 2581 1326
rect 2594 1293 2597 1326
rect 2626 1313 2629 1426
rect 2546 1103 2549 1196
rect 2562 1193 2565 1216
rect 2594 1196 2597 1206
rect 2570 1143 2573 1156
rect 2554 1113 2557 1126
rect 2562 1123 2573 1126
rect 2562 1113 2565 1123
rect 2578 1076 2581 1196
rect 2594 1193 2613 1196
rect 2570 1073 2581 1076
rect 2506 1013 2509 1036
rect 2498 903 2501 1006
rect 2498 733 2501 886
rect 2506 776 2509 986
rect 2514 963 2517 1016
rect 2514 893 2517 926
rect 2522 883 2525 1016
rect 2538 993 2541 1006
rect 2562 996 2565 1036
rect 2570 1006 2573 1073
rect 2586 1066 2589 1136
rect 2578 1063 2589 1066
rect 2578 1033 2581 1063
rect 2594 1056 2597 1126
rect 2602 1103 2605 1116
rect 2610 1103 2613 1193
rect 2618 1136 2621 1216
rect 2626 1143 2637 1146
rect 2618 1133 2629 1136
rect 2618 1113 2621 1126
rect 2586 1053 2597 1056
rect 2578 1013 2581 1026
rect 2570 1003 2581 1006
rect 2586 1003 2589 1053
rect 2594 1013 2597 1036
rect 2554 986 2557 996
rect 2562 993 2573 996
rect 2554 983 2565 986
rect 2538 933 2541 966
rect 2530 863 2533 916
rect 2506 773 2533 776
rect 2530 733 2533 773
rect 2538 753 2541 926
rect 2546 896 2549 936
rect 2554 923 2557 976
rect 2562 933 2565 983
rect 2570 933 2573 993
rect 2578 933 2581 1003
rect 2602 963 2605 1006
rect 2594 933 2605 936
rect 2578 903 2581 916
rect 2546 893 2557 896
rect 2554 846 2557 893
rect 2594 866 2597 926
rect 2546 843 2557 846
rect 2586 863 2597 866
rect 2546 793 2549 843
rect 2562 823 2581 826
rect 2562 813 2565 823
rect 2578 733 2581 816
rect 2586 813 2589 863
rect 2602 826 2605 926
rect 2594 823 2605 826
rect 2594 813 2597 823
rect 2586 793 2589 806
rect 2602 743 2605 816
rect 2610 813 2613 1096
rect 2618 1083 2621 1106
rect 2618 983 2621 1016
rect 2626 1003 2629 1133
rect 2634 1113 2637 1136
rect 2642 1093 2645 1516
rect 2658 1496 2661 1586
rect 2654 1493 2661 1496
rect 2654 1216 2657 1493
rect 2654 1213 2661 1216
rect 2650 1076 2653 1196
rect 2642 1073 2653 1076
rect 2642 1003 2645 1073
rect 2658 1056 2661 1213
rect 2654 1053 2661 1056
rect 2654 966 2657 1053
rect 2654 963 2661 966
rect 2634 923 2645 926
rect 2658 813 2661 963
rect 2610 793 2613 806
rect 2434 713 2445 716
rect 2466 713 2469 726
rect 2498 723 2509 726
rect 2514 723 2533 726
rect 2498 646 2501 723
rect 2514 716 2517 723
rect 2466 633 2469 646
rect 2490 643 2501 646
rect 2506 713 2517 716
rect 2442 546 2445 606
rect 2402 543 2421 546
rect 2434 543 2445 546
rect 2402 533 2405 543
rect 2410 433 2413 446
rect 2402 423 2413 426
rect 2418 416 2421 526
rect 2434 493 2437 543
rect 2450 536 2453 626
rect 2442 533 2453 536
rect 2458 516 2461 616
rect 2482 583 2485 636
rect 2490 603 2493 643
rect 2498 623 2501 636
rect 2506 606 2509 713
rect 2514 693 2517 706
rect 2522 633 2525 716
rect 2586 693 2589 736
rect 2594 733 2605 736
rect 2666 733 2669 1593
rect 2522 623 2541 626
rect 2522 613 2525 623
rect 2538 616 2541 623
rect 2562 616 2565 626
rect 2538 613 2549 616
rect 2554 613 2565 616
rect 2450 513 2461 516
rect 2466 523 2493 526
rect 2498 523 2501 606
rect 2506 603 2525 606
rect 2506 533 2509 546
rect 2450 446 2453 513
rect 2450 443 2461 446
rect 2426 423 2429 436
rect 2410 413 2421 416
rect 2402 316 2405 386
rect 2410 333 2413 356
rect 2434 323 2437 436
rect 2442 413 2445 426
rect 2450 406 2453 426
rect 2458 423 2461 443
rect 2466 413 2469 523
rect 2474 423 2477 516
rect 2490 436 2493 506
rect 2498 503 2501 516
rect 2506 476 2509 526
rect 2514 493 2517 603
rect 2530 593 2533 606
rect 2538 603 2549 606
rect 2522 543 2525 586
rect 2522 503 2525 526
rect 2538 486 2541 526
rect 2530 483 2541 486
rect 2506 473 2517 476
rect 2490 433 2501 436
rect 2450 403 2461 406
rect 2482 403 2485 416
rect 2490 403 2493 433
rect 2498 403 2501 416
rect 2506 403 2509 416
rect 2514 396 2517 473
rect 2530 436 2533 483
rect 2530 433 2541 436
rect 2538 413 2541 433
rect 2546 413 2549 596
rect 2554 423 2557 613
rect 2562 593 2565 606
rect 2570 576 2573 606
rect 2578 603 2581 616
rect 2594 613 2597 646
rect 2586 603 2597 606
rect 2562 573 2573 576
rect 2562 533 2565 573
rect 2578 543 2581 586
rect 2570 523 2573 536
rect 2586 526 2589 603
rect 2582 523 2589 526
rect 2582 456 2585 523
rect 2582 453 2589 456
rect 2562 423 2565 436
rect 2570 426 2573 446
rect 2586 436 2589 453
rect 2578 433 2589 436
rect 2570 423 2581 426
rect 2506 393 2525 396
rect 2442 333 2445 346
rect 2450 333 2453 366
rect 2522 356 2525 393
rect 2522 353 2533 356
rect 2402 313 2413 316
rect 2386 303 2405 306
rect 2354 233 2365 236
rect 2410 233 2413 313
rect 2306 193 2309 206
rect 2338 203 2341 216
rect 2314 193 2325 196
rect 2314 163 2317 193
rect 2330 183 2333 196
rect 2354 193 2357 233
rect 2362 203 2365 216
rect 2370 213 2373 226
rect 2402 213 2405 226
rect 2418 203 2421 306
rect 2426 303 2429 316
rect 2466 246 2469 336
rect 2482 323 2485 336
rect 2490 323 2509 326
rect 2474 313 2485 316
rect 2482 246 2485 313
rect 2490 303 2493 316
rect 2514 256 2517 336
rect 2522 333 2525 353
rect 2538 313 2541 406
rect 2554 323 2557 416
rect 2562 413 2573 416
rect 2570 333 2573 346
rect 2578 323 2581 423
rect 2586 316 2589 426
rect 2594 403 2597 596
rect 2602 593 2605 726
rect 2618 696 2621 726
rect 2614 693 2621 696
rect 2614 616 2617 693
rect 2610 613 2617 616
rect 2610 583 2613 613
rect 2618 593 2621 606
rect 2626 603 2629 726
rect 2634 613 2637 626
rect 2610 466 2613 526
rect 2642 523 2645 616
rect 2610 463 2621 466
rect 2594 333 2597 356
rect 2602 333 2605 436
rect 2618 403 2621 463
rect 2626 403 2629 456
rect 2650 356 2653 426
rect 2650 353 2661 356
rect 2658 333 2661 353
rect 2570 313 2589 316
rect 2506 253 2517 256
rect 2466 243 2477 246
rect 2482 243 2493 246
rect 2426 193 2429 236
rect 2434 213 2437 226
rect 2442 206 2445 216
rect 2434 203 2445 206
rect 2434 173 2437 203
rect 2442 183 2445 196
rect 2458 193 2461 206
rect 2474 196 2477 243
rect 2490 216 2493 243
rect 2490 213 2501 216
rect 2506 213 2509 253
rect 2514 213 2517 226
rect 2538 213 2541 226
rect 2546 223 2549 306
rect 2546 213 2565 216
rect 2498 206 2501 213
rect 2482 203 2493 206
rect 2498 203 2517 206
rect 2474 193 2485 196
rect 2538 183 2541 206
rect 2578 193 2581 206
rect 2626 193 2629 206
rect 2290 73 2293 116
rect 690 13 701 16
rect 690 -88 693 13
rect 1224 -19 1227 38
rect 2678 37 2698 2603
rect 2702 13 2722 2627
rect 2730 1533 2733 2136
rect 2742 1040 2745 2637
rect 2749 1340 2752 2645
rect 2756 1641 2759 2653
rect 2764 1941 2767 2661
rect 2774 2240 2777 2670
rect 2785 2540 2788 2683
rect 2785 2537 2859 2540
rect 2848 2473 2858 2476
rect 2774 2237 2859 2240
rect 2848 2173 2859 2176
rect 2764 1938 2860 1941
rect 2848 1872 2858 1875
rect 2756 1638 2859 1641
rect 2848 1572 2859 1575
rect 2749 1337 2859 1340
rect 2848 1273 2859 1276
rect 2742 1037 2859 1040
rect 2849 673 2859 676
rect 2800 649 2860 652
rect 2800 -88 2803 649
rect 2849 372 2858 375
rect 690 -91 2803 -88
rect 2810 349 2859 352
rect 2810 -96 2813 349
rect 2849 72 2859 75
rect 674 -99 2813 -96
rect 2823 51 2860 54
rect 2823 -106 2826 51
rect 658 -109 2826 -106
rect 642 -119 1074 -116
rect 474 -128 1067 -125
rect 458 -138 1061 -135
rect 290 -144 1055 -141
rect 202 -150 1049 -147
rect -68 -156 525 -153
rect -74 -162 226 -159
rect 199 -184 202 -175
rect 223 -185 226 -162
rect 500 -184 503 -175
rect 522 -184 525 -156
rect 1046 -158 1049 -150
rect 1052 -151 1055 -144
rect 1058 -145 1061 -138
rect 1064 -137 1067 -128
rect 1071 -131 1074 -119
rect 1071 -134 1453 -131
rect 1064 -140 1446 -137
rect 1058 -148 1438 -145
rect 1052 -154 1432 -151
rect 1429 -158 1432 -154
rect 1435 -152 1438 -148
rect 1443 -146 1446 -140
rect 1450 -140 1453 -134
rect 1450 -143 1743 -140
rect 1740 -145 1743 -143
rect 1443 -149 1737 -146
rect 1740 -148 2039 -145
rect 1734 -152 1737 -149
rect 2036 -151 2039 -148
rect 1435 -155 1731 -152
rect 1734 -155 2032 -152
rect 2036 -154 2332 -151
rect 1728 -158 1731 -155
rect 2029 -158 2032 -155
rect 2329 -158 2332 -154
rect 1046 -161 1426 -158
rect 1429 -161 1725 -158
rect 1728 -161 2025 -158
rect 2029 -161 2325 -158
rect 2329 -161 2627 -158
rect 799 -184 802 -175
rect 1035 -184 1038 -162
rect 1399 -184 1402 -174
rect 1423 -184 1426 -161
rect 1699 -184 1702 -174
rect 1722 -184 1725 -161
rect 1999 -184 2002 -174
rect 2022 -184 2025 -161
rect 2299 -184 2302 -174
rect 2322 -184 2325 -161
rect 2599 -184 2602 -174
rect 2624 -185 2627 -161
<< m3contact >>
rect 433 2741 438 2746
rect 733 2739 738 2744
rect 1034 2741 1039 2746
rect 1111 2742 1116 2747
rect -38 2536 -33 2541
rect -18 2651 -13 2656
rect -8 2643 -3 2648
rect 0 2402 5 2407
rect -7 2202 -2 2207
rect -8 2182 -3 2187
rect 0 2132 5 2137
rect -26 1269 -21 1274
rect 0 1322 5 1327
rect 0 1268 5 1273
rect -12 1142 -7 1147
rect 0 1002 5 1007
rect 0 812 5 817
rect 0 732 5 737
rect 0 712 5 717
rect -88 637 -83 642
rect 0 532 5 537
rect -88 335 -83 340
rect 0 332 5 337
rect 0 172 5 177
rect 1035 -162 1040 -157
<< metal3 >>
rect 1110 2747 1117 2748
rect 432 2746 439 2747
rect 432 2741 433 2746
rect 438 2741 439 2746
rect 1033 2746 1040 2747
rect 432 2740 439 2741
rect 732 2744 739 2745
rect 433 2665 438 2740
rect 732 2739 733 2744
rect 738 2739 739 2744
rect 1033 2741 1034 2746
rect 1039 2741 1040 2746
rect 1110 2742 1111 2747
rect 1116 2742 1117 2747
rect 1110 2741 1117 2742
rect 1033 2740 1040 2741
rect 732 2738 739 2739
rect -27 2660 438 2665
rect -27 2647 -22 2660
rect 733 2657 738 2738
rect -19 2656 738 2657
rect -19 2651 -18 2656
rect -13 2652 738 2656
rect -13 2651 -12 2652
rect -19 2650 -12 2651
rect 1034 2649 1039 2740
rect -9 2648 1039 2649
rect -27 2642 -14 2647
rect -9 2643 -8 2648
rect -3 2644 1039 2648
rect -3 2643 -2 2644
rect -9 2642 -2 2643
rect -39 2541 -32 2542
rect -39 2536 -38 2541
rect -33 2536 -23 2541
rect -39 2535 -32 2536
rect -28 2117 -23 2536
rect -19 2157 -14 2642
rect 1111 2639 1116 2741
rect -11 2634 1116 2639
rect -11 2337 -6 2634
rect 801 2602 1110 2607
rect 801 2597 806 2602
rect 577 2592 806 2597
rect 577 2587 582 2592
rect 1105 2587 1110 2602
rect 561 2582 582 2587
rect 841 2582 1070 2587
rect 1105 2582 1334 2587
rect 561 2572 566 2582
rect 841 2577 846 2582
rect 817 2572 846 2577
rect 1065 2577 1070 2582
rect 1065 2572 1094 2577
rect 593 2562 990 2567
rect 1041 2562 1078 2567
rect 1873 2562 2046 2567
rect 593 2557 598 2562
rect 577 2552 598 2557
rect 801 2552 854 2557
rect 1089 2552 1166 2557
rect 1321 2552 1350 2557
rect 1377 2552 1446 2557
rect 1505 2552 1694 2557
rect 177 2542 486 2547
rect 625 2542 686 2547
rect 713 2542 822 2547
rect 841 2542 886 2547
rect 1033 2542 1118 2547
rect 1193 2542 1254 2547
rect 1305 2542 1494 2547
rect 1505 2537 1510 2552
rect 1689 2547 1694 2552
rect 1873 2547 1878 2562
rect 1689 2542 1718 2547
rect 1849 2542 1878 2547
rect 2041 2547 2046 2562
rect 2401 2552 2454 2557
rect 2041 2542 2102 2547
rect 2249 2542 2502 2547
rect 449 2532 614 2537
rect 705 2532 1510 2537
rect 1825 2532 2030 2537
rect 2281 2532 2310 2537
rect 2345 2532 2550 2537
rect 609 2527 710 2532
rect 729 2522 862 2527
rect 1081 2522 1606 2527
rect 1617 2522 1726 2527
rect 1881 2522 1982 2527
rect 2297 2522 2374 2527
rect 2425 2522 2470 2527
rect 2481 2522 2486 2532
rect 2505 2522 2566 2527
rect 1617 2517 1622 2522
rect 225 2512 278 2517
rect 665 2512 790 2517
rect 873 2512 1070 2517
rect 1329 2512 1382 2517
rect 1409 2512 1622 2517
rect 1633 2512 1726 2517
rect 1777 2512 1870 2517
rect 2129 2512 2246 2517
rect 2361 2512 2430 2517
rect 2441 2512 2542 2517
rect 785 2507 878 2512
rect 1065 2507 1334 2512
rect 2129 2507 2134 2512
rect 497 2502 646 2507
rect 721 2502 766 2507
rect 1353 2502 1382 2507
rect 1553 2502 2134 2507
rect 2241 2507 2246 2512
rect 2241 2502 2422 2507
rect 2473 2502 2510 2507
rect 497 2497 502 2502
rect 473 2492 502 2497
rect 641 2497 646 2502
rect 1377 2497 1558 2502
rect 641 2492 1206 2497
rect 1225 2492 1334 2497
rect 1577 2492 1606 2497
rect 1225 2487 1230 2492
rect 353 2482 630 2487
rect 1121 2482 1230 2487
rect 1329 2487 1334 2492
rect 1601 2487 1606 2492
rect 1665 2492 1702 2497
rect 1769 2492 1934 2497
rect 2169 2492 2198 2497
rect 1665 2487 1670 2492
rect 2193 2487 2198 2492
rect 2329 2492 2438 2497
rect 2329 2487 2334 2492
rect 1329 2482 1390 2487
rect 1409 2482 1534 2487
rect 1601 2482 1670 2487
rect 1689 2482 1758 2487
rect 1945 2482 2038 2487
rect 625 2477 630 2482
rect 913 2477 1126 2482
rect 1409 2477 1414 2482
rect 465 2472 494 2477
rect 625 2472 918 2477
rect 1145 2472 1414 2477
rect 1529 2477 1534 2482
rect 1753 2477 1950 2482
rect 2033 2477 2038 2482
rect 2145 2482 2174 2487
rect 2193 2482 2334 2487
rect 2145 2477 2150 2482
rect 1529 2472 1558 2477
rect 2033 2472 2150 2477
rect 937 2462 1046 2467
rect 1041 2457 1046 2462
rect 1169 2462 1662 2467
rect 1777 2462 1942 2467
rect 1169 2457 1174 2462
rect 609 2452 694 2457
rect 825 2452 878 2457
rect 905 2452 942 2457
rect 1041 2452 1174 2457
rect 1249 2452 1302 2457
rect 1425 2452 1822 2457
rect 1921 2452 2014 2457
rect 2489 2452 2534 2457
rect 609 2447 614 2452
rect 497 2442 614 2447
rect 689 2447 694 2452
rect 1297 2447 1430 2452
rect 689 2442 718 2447
rect 841 2442 902 2447
rect 969 2442 1022 2447
rect 1193 2442 1278 2447
rect 1449 2442 1606 2447
rect 1809 2442 1966 2447
rect 1977 2442 2046 2447
rect 1369 2432 1446 2437
rect 1809 2432 1846 2437
rect 1929 2432 2022 2437
rect 2033 2432 2166 2437
rect 2281 2432 2318 2437
rect 2601 2432 2662 2437
rect 1441 2427 1446 2432
rect 97 2422 198 2427
rect 209 2422 518 2427
rect 625 2422 790 2427
rect 801 2422 838 2427
rect 953 2422 1014 2427
rect 1161 2422 1422 2427
rect 1441 2422 1558 2427
rect 1569 2422 1622 2427
rect 1641 2422 1678 2427
rect 1705 2422 1758 2427
rect 1785 2422 1822 2427
rect 1937 2422 1998 2427
rect 2337 2422 2414 2427
rect 2497 2422 2550 2427
rect 1553 2417 1558 2422
rect 2017 2417 2110 2422
rect 2337 2417 2342 2422
rect 585 2412 638 2417
rect 681 2412 734 2417
rect 921 2412 950 2417
rect 1049 2412 1078 2417
rect 1201 2412 1326 2417
rect 1553 2412 1670 2417
rect -1 2407 6 2408
rect 105 2407 262 2412
rect 945 2407 1054 2412
rect -1 2402 0 2407
rect 5 2402 70 2407
rect 81 2402 110 2407
rect 257 2402 286 2407
rect 305 2402 502 2407
rect 697 2402 838 2407
rect 1121 2402 1182 2407
rect -1 2401 6 2402
rect 65 2392 70 2402
rect 145 2392 222 2397
rect 545 2392 630 2397
rect 641 2392 758 2397
rect 833 2392 838 2402
rect 1665 2397 1670 2412
rect 1833 2412 2022 2417
rect 2105 2412 2134 2417
rect 2177 2412 2342 2417
rect 2409 2417 2414 2422
rect 2409 2412 2518 2417
rect 2561 2412 2582 2417
rect 1833 2397 1838 2412
rect 2129 2407 2134 2412
rect 1889 2402 2118 2407
rect 2129 2402 2150 2407
rect 2145 2397 2150 2402
rect 2225 2402 2254 2407
rect 2497 2402 2574 2407
rect 2225 2397 2230 2402
rect 969 2392 1038 2397
rect 1433 2392 1518 2397
rect 1665 2392 1838 2397
rect 1937 2392 1990 2397
rect 2145 2392 2230 2397
rect 2337 2392 2454 2397
rect 2497 2392 2622 2397
rect 1433 2387 1438 2392
rect 241 2382 374 2387
rect 561 2382 742 2387
rect 761 2382 846 2387
rect 865 2382 942 2387
rect 1001 2382 1046 2387
rect 1065 2382 1142 2387
rect 1337 2382 1438 2387
rect 1513 2387 1518 2392
rect 2497 2387 2502 2392
rect 1513 2382 1638 2387
rect 2017 2382 2118 2387
rect 2369 2382 2502 2387
rect 2521 2382 2542 2387
rect 241 2377 246 2382
rect 185 2372 246 2377
rect 369 2377 374 2382
rect 1065 2377 1070 2382
rect 369 2372 550 2377
rect 649 2372 718 2377
rect 1009 2372 1070 2377
rect 1137 2377 1142 2382
rect 1137 2372 1166 2377
rect 1281 2372 1334 2377
rect 1425 2372 1502 2377
rect 1617 2372 1646 2377
rect 1857 2372 1926 2377
rect 81 2362 358 2367
rect 545 2357 550 2372
rect 865 2367 990 2372
rect 1921 2367 1926 2372
rect 2001 2372 2030 2377
rect 2241 2372 2350 2377
rect 2481 2372 2566 2377
rect 2001 2367 2006 2372
rect 609 2362 758 2367
rect 769 2362 806 2367
rect 841 2362 870 2367
rect 985 2362 1350 2367
rect 1737 2362 1838 2367
rect 1921 2362 2006 2367
rect 2169 2362 2342 2367
rect 2433 2362 2478 2367
rect 161 2352 238 2357
rect 369 2352 526 2357
rect 545 2352 1222 2357
rect 1697 2352 1766 2357
rect 2201 2352 2238 2357
rect 65 2337 70 2347
rect 145 2342 222 2347
rect 337 2342 398 2347
rect 473 2342 550 2347
rect 1313 2342 1358 2347
rect 1481 2342 1558 2347
rect 1801 2342 1822 2347
rect 569 2337 814 2342
rect 873 2337 990 2342
rect 1065 2337 1294 2342
rect -11 2332 70 2337
rect 81 2332 110 2337
rect 105 2317 110 2332
rect 233 2332 302 2337
rect 465 2332 574 2337
rect 809 2332 878 2337
rect 985 2332 1014 2337
rect 1041 2332 1070 2337
rect 1289 2332 1470 2337
rect 1537 2332 1566 2337
rect 1729 2332 1750 2337
rect 1929 2332 2046 2337
rect 2161 2332 2238 2337
rect 233 2317 238 2332
rect 1465 2327 1542 2332
rect 2161 2327 2166 2332
rect 505 2322 798 2327
rect 889 2322 966 2327
rect 1089 2322 1422 2327
rect 1585 2322 1710 2327
rect 1881 2322 1918 2327
rect 1953 2322 2166 2327
rect 2233 2327 2238 2332
rect 2489 2332 2566 2337
rect 2489 2327 2494 2332
rect 2233 2322 2262 2327
rect 2273 2322 2366 2327
rect 2465 2322 2494 2327
rect 2561 2327 2566 2332
rect 2561 2322 2590 2327
rect 793 2317 894 2322
rect 961 2317 1094 2322
rect 1585 2317 1590 2322
rect 1705 2317 1790 2322
rect 105 2312 238 2317
rect 345 2312 470 2317
rect 713 2312 774 2317
rect 913 2312 942 2317
rect 937 2307 942 2312
rect 1113 2312 1190 2317
rect 1369 2312 1422 2317
rect 1441 2312 1590 2317
rect 1785 2312 1870 2317
rect 1113 2307 1118 2312
rect 1185 2307 1374 2312
rect 1865 2307 1870 2312
rect 1953 2307 1958 2322
rect 1977 2312 2078 2317
rect 2177 2312 2246 2317
rect 2273 2312 2278 2322
rect 2297 2312 2518 2317
rect 489 2302 518 2307
rect 665 2302 766 2307
rect 785 2302 838 2307
rect 857 2302 902 2307
rect 937 2302 1118 2307
rect 1137 2302 1166 2307
rect 1161 2297 1166 2302
rect 1393 2302 1470 2307
rect 1593 2302 1638 2307
rect 1665 2302 1774 2307
rect 1865 2302 1958 2307
rect 2209 2302 2438 2307
rect 2521 2302 2558 2307
rect 1393 2297 1398 2302
rect 537 2292 646 2297
rect 745 2292 790 2297
rect 865 2292 910 2297
rect 1161 2292 1398 2297
rect 1609 2292 1638 2297
rect 1753 2292 1782 2297
rect 2185 2292 2214 2297
rect 537 2287 542 2292
rect 337 2282 542 2287
rect 641 2287 646 2292
rect 1441 2287 1590 2292
rect 1633 2287 1758 2292
rect 2209 2287 2214 2292
rect 2337 2292 2366 2297
rect 2417 2292 2454 2297
rect 2337 2287 2342 2292
rect 641 2282 846 2287
rect 929 2282 1118 2287
rect 1417 2282 1446 2287
rect 1585 2282 1614 2287
rect 249 2272 430 2277
rect 777 2272 806 2277
rect 929 2272 934 2282
rect 1113 2277 1118 2282
rect 1609 2277 1614 2282
rect 1793 2282 2070 2287
rect 2209 2282 2342 2287
rect 1793 2277 1798 2282
rect 1113 2272 1398 2277
rect 833 2267 934 2272
rect 1393 2267 1398 2272
rect 1457 2272 1590 2277
rect 1609 2272 1798 2277
rect 1457 2267 1462 2272
rect 185 2262 374 2267
rect 369 2257 374 2262
rect 441 2262 486 2267
rect 441 2257 446 2262
rect 369 2252 446 2257
rect 481 2247 486 2262
rect 601 2262 838 2267
rect 1393 2262 1462 2267
rect 1473 2262 1566 2267
rect 601 2247 606 2262
rect 697 2252 726 2257
rect 817 2252 846 2257
rect 889 2252 1382 2257
rect 1577 2252 1950 2257
rect 721 2247 822 2252
rect 1377 2247 1582 2252
rect 257 2242 350 2247
rect 481 2242 606 2247
rect 625 2242 702 2247
rect 2209 2242 2366 2247
rect 2449 2242 2510 2247
rect 1041 2237 1358 2242
rect 281 2232 462 2237
rect 625 2232 830 2237
rect 929 2232 1046 2237
rect 1353 2232 1446 2237
rect 1537 2232 1590 2237
rect 2353 2232 2390 2237
rect 2473 2232 2590 2237
rect 1441 2227 1446 2232
rect 105 2222 238 2227
rect 313 2222 366 2227
rect 377 2222 406 2227
rect 401 2217 406 2222
rect 473 2222 534 2227
rect 633 2222 678 2227
rect 1057 2222 1342 2227
rect 1441 2222 1878 2227
rect 473 2217 478 2222
rect 241 2212 374 2217
rect 401 2212 478 2217
rect 809 2212 846 2217
rect 929 2212 1150 2217
rect 1233 2212 1310 2217
rect 1785 2212 1806 2217
rect -8 2207 -1 2208
rect 153 2207 222 2212
rect 1497 2207 1590 2212
rect -8 2202 -7 2207
rect -2 2202 158 2207
rect 217 2202 262 2207
rect -8 2201 -1 2202
rect 169 2192 230 2197
rect 257 2192 262 2202
rect 561 2202 1142 2207
rect 1185 2202 1214 2207
rect 1313 2202 1366 2207
rect 1473 2202 1502 2207
rect 1585 2202 1670 2207
rect 1713 2202 1862 2207
rect 561 2197 566 2202
rect 1185 2197 1190 2202
rect 1473 2197 1478 2202
rect 345 2192 566 2197
rect 577 2192 606 2197
rect 769 2192 814 2197
rect -9 2187 -2 2188
rect 625 2187 734 2192
rect 809 2187 814 2192
rect 953 2192 982 2197
rect 1009 2192 1030 2197
rect 1041 2192 1086 2197
rect 1169 2192 1190 2197
rect 1209 2192 1478 2197
rect 1497 2192 1574 2197
rect 1641 2192 1750 2197
rect 1761 2192 1870 2197
rect 953 2187 958 2192
rect -9 2182 -8 2187
rect -3 2182 70 2187
rect 257 2182 630 2187
rect 729 2182 790 2187
rect 809 2182 958 2187
rect 1025 2187 1030 2192
rect 1025 2182 1302 2187
rect -9 2181 -2 2182
rect 1297 2177 1302 2182
rect 1473 2182 1894 2187
rect 1905 2182 1910 2227
rect 1921 2182 1926 2227
rect 1969 2207 1974 2227
rect 1953 2202 1974 2207
rect 1953 2187 1958 2202
rect 1953 2182 1982 2187
rect 2097 2182 2102 2227
rect 2353 2222 2462 2227
rect 2273 2207 2278 2217
rect 2369 2212 2398 2217
rect 2241 2202 2278 2207
rect 2393 2207 2398 2212
rect 2473 2212 2502 2217
rect 2473 2207 2478 2212
rect 2393 2202 2478 2207
rect 2225 2192 2326 2197
rect 2185 2182 2294 2187
rect 2561 2182 2566 2227
rect 1473 2177 1478 2182
rect 113 2172 254 2177
rect 393 2172 454 2177
rect 617 2172 718 2177
rect 1145 2172 1278 2177
rect 1297 2172 1478 2177
rect 1529 2172 1766 2177
rect 1873 2172 2046 2177
rect 977 2167 1078 2172
rect 161 2157 262 2162
rect 433 2157 438 2167
rect 449 2162 630 2167
rect 673 2162 982 2167
rect 1073 2162 1142 2167
rect 1497 2162 1614 2167
rect 1665 2162 1918 2167
rect 1137 2157 1142 2162
rect -19 2152 166 2157
rect 257 2152 286 2157
rect 433 2152 462 2157
rect 609 2152 646 2157
rect 657 2152 694 2157
rect 993 2152 1062 2157
rect 1137 2152 1286 2157
rect 1329 2152 1422 2157
rect 1505 2152 1654 2157
rect 1665 2152 1694 2157
rect 1753 2152 1814 2157
rect 1825 2152 1894 2157
rect 1913 2147 1918 2162
rect 2057 2162 2182 2167
rect 2513 2162 2614 2167
rect 2057 2147 2062 2162
rect 2281 2152 2334 2157
rect 2369 2152 2486 2157
rect 2593 2152 2630 2157
rect 2369 2147 2374 2152
rect 177 2142 238 2147
rect 321 2142 350 2147
rect 1481 2142 1574 2147
rect 1641 2142 1678 2147
rect 1745 2142 1846 2147
rect 1913 2142 2062 2147
rect 2129 2142 2150 2147
rect 2257 2142 2374 2147
rect -1 2137 6 2138
rect 233 2137 326 2142
rect -1 2132 0 2137
rect 5 2132 94 2137
rect 409 2132 454 2137
rect 521 2132 566 2137
rect 697 2132 742 2137
rect -1 2131 6 2132
rect 137 2122 198 2127
rect 233 2122 262 2127
rect 585 2122 646 2127
rect 681 2122 702 2127
rect 737 2122 742 2132
rect 809 2132 974 2137
rect 1041 2132 1078 2137
rect 809 2127 814 2132
rect 785 2122 814 2127
rect 969 2127 974 2132
rect 1537 2127 1542 2137
rect 1689 2132 1838 2137
rect 969 2122 1206 2127
rect 1225 2122 1462 2127
rect 1537 2122 1598 2127
rect 1777 2122 1822 2127
rect 2129 2122 2134 2142
rect 2233 2132 2310 2137
rect 2321 2132 2382 2137
rect 2289 2122 2358 2127
rect 2385 2122 2414 2127
rect 1225 2117 1230 2122
rect -28 2112 70 2117
rect 209 2112 486 2117
rect 625 2112 678 2117
rect 689 2112 718 2117
rect 1041 2112 1230 2117
rect 1457 2107 1462 2122
rect 2497 2117 2502 2147
rect 2625 2137 2630 2152
rect 2625 2132 2662 2137
rect 1481 2112 1518 2117
rect 1529 2112 1574 2117
rect 1633 2112 1670 2117
rect 1761 2112 1830 2117
rect 1897 2112 2110 2117
rect 2145 2112 2174 2117
rect 2465 2112 2502 2117
rect 2601 2112 2670 2117
rect 233 2102 294 2107
rect 353 2102 382 2107
rect 497 2102 1014 2107
rect 377 2097 502 2102
rect 1009 2097 1014 2102
rect 1113 2102 1398 2107
rect 1457 2102 1558 2107
rect 1705 2102 1878 2107
rect 1113 2097 1118 2102
rect 1553 2097 1686 2102
rect 1897 2097 1902 2112
rect 649 2092 686 2097
rect 1009 2092 1118 2097
rect 1185 2092 1246 2097
rect 1273 2092 1310 2097
rect 1465 2092 1542 2097
rect 1681 2092 1902 2097
rect 2105 2097 2110 2112
rect 2193 2102 2278 2107
rect 2321 2102 2406 2107
rect 2273 2097 2278 2102
rect 2105 2092 2214 2097
rect 2273 2092 2318 2097
rect 553 2087 630 2092
rect 305 2082 374 2087
rect 489 2082 558 2087
rect 625 2082 798 2087
rect 1137 2082 1214 2087
rect 1417 2082 2286 2087
rect 569 2072 654 2077
rect 817 2072 990 2077
rect 1361 2072 1614 2077
rect 1745 2072 1942 2077
rect 761 2062 790 2067
rect 585 2057 678 2062
rect 817 2057 822 2072
rect 985 2057 990 2072
rect 1609 2067 1750 2072
rect 1089 2062 1222 2067
rect 1417 2062 1590 2067
rect 1585 2057 1590 2062
rect 1769 2062 1798 2067
rect 1873 2062 1910 2067
rect 1769 2057 1774 2062
rect 561 2052 590 2057
rect 673 2052 822 2057
rect 841 2052 910 2057
rect 985 2052 1118 2057
rect 1257 2052 1342 2057
rect 1441 2052 1494 2057
rect 1521 2052 1566 2057
rect 1585 2052 1774 2057
rect 1937 2057 1942 2072
rect 2097 2072 2190 2077
rect 2097 2057 2102 2072
rect 1937 2052 2102 2057
rect 2457 2052 2550 2057
rect 841 2047 846 2052
rect 273 2042 366 2047
rect 625 2042 662 2047
rect 753 2042 846 2047
rect 905 2047 910 2052
rect 2457 2047 2462 2052
rect 905 2042 998 2047
rect 1153 2042 1190 2047
rect 1297 2042 1414 2047
rect 1449 2042 1566 2047
rect 2121 2042 2166 2047
rect 2433 2042 2462 2047
rect 2545 2047 2550 2052
rect 2545 2042 2582 2047
rect 657 2037 758 2042
rect 1153 2037 1158 2042
rect 1409 2037 1414 2042
rect 425 2032 638 2037
rect 777 2032 894 2037
rect 969 2032 1158 2037
rect 1177 2032 1302 2037
rect 1337 2032 1398 2037
rect 1409 2032 1478 2037
rect 1489 2032 1518 2037
rect 1585 2032 1614 2037
rect 1649 2032 1710 2037
rect 1777 2032 1918 2037
rect 2361 2032 2446 2037
rect 617 2012 678 2017
rect 441 2002 470 2007
rect 481 2002 542 2007
rect 593 2002 694 2007
rect 737 1997 742 2027
rect 785 2022 814 2027
rect 1105 2022 1190 2027
rect 1305 2022 1430 2027
rect 833 2017 958 2022
rect 769 2012 838 2017
rect 953 2012 982 2017
rect 1073 2012 1158 2017
rect 793 2002 862 2007
rect 889 2002 1062 2007
rect 1169 2002 1310 2007
rect 1057 1997 1174 2002
rect 241 1992 358 1997
rect 369 1992 518 1997
rect 577 1992 686 1997
rect 737 1992 798 1997
rect 953 1992 998 1997
rect 1393 1987 1398 2017
rect 1441 2007 1446 2027
rect 1457 2022 1478 2027
rect 1497 2022 1582 2027
rect 1881 2022 1926 2027
rect 2009 2022 2158 2027
rect 2185 2022 2230 2027
rect 2297 2022 2382 2027
rect 2465 2022 2502 2027
rect 1473 2017 1478 2022
rect 1473 2012 1646 2017
rect 1793 2012 1870 2017
rect 1441 2002 1518 2007
rect 1537 2002 1638 2007
rect 1817 2002 1894 2007
rect 2497 1992 2502 2022
rect 209 1982 270 1987
rect 449 1982 518 1987
rect 593 1982 910 1987
rect 977 1982 1310 1987
rect 1353 1982 1558 1987
rect 1569 1982 1630 1987
rect 1721 1982 1806 1987
rect 1977 1982 2030 1987
rect 2161 1982 2254 1987
rect 2321 1982 2358 1987
rect 2529 1982 2534 2027
rect 2641 2022 2662 2027
rect 2609 2012 2638 2017
rect 2657 2002 2662 2022
rect 593 1977 598 1982
rect 1553 1977 1558 1982
rect 161 1972 374 1977
rect 489 1972 598 1977
rect 609 1972 710 1977
rect 753 1972 782 1977
rect 817 1972 886 1977
rect 1217 1972 1286 1977
rect 1553 1972 1742 1977
rect 1841 1972 1910 1977
rect 2217 1972 2286 1977
rect 1217 1967 1222 1972
rect 1281 1967 1430 1972
rect 377 1962 406 1967
rect 457 1962 718 1967
rect 761 1962 814 1967
rect 1009 1962 1038 1967
rect 1105 1962 1222 1967
rect 1233 1962 1270 1967
rect 1425 1962 1542 1967
rect 1617 1962 1646 1967
rect 1929 1962 1958 1967
rect 2129 1962 2174 1967
rect 1537 1957 1622 1962
rect 73 1952 246 1957
rect 345 1952 398 1957
rect 513 1952 574 1957
rect 641 1952 702 1957
rect 761 1952 1102 1957
rect 1185 1952 1262 1957
rect 1297 1952 1414 1957
rect 1681 1952 1838 1957
rect 1881 1952 1918 1957
rect 1681 1947 1686 1952
rect 185 1942 230 1947
rect 313 1942 406 1947
rect 553 1942 614 1947
rect 633 1942 758 1947
rect 833 1942 902 1947
rect 961 1942 1030 1947
rect 1089 1942 1174 1947
rect 1505 1942 1686 1947
rect 1833 1947 1838 1952
rect 1937 1947 1942 1957
rect 1833 1942 1942 1947
rect 129 1932 310 1937
rect 121 1922 174 1927
rect 225 1922 254 1927
rect 305 1922 310 1932
rect 361 1922 382 1927
rect 233 1912 286 1917
rect 297 1912 334 1917
rect 401 1912 406 1942
rect 753 1937 758 1942
rect 1169 1937 1278 1942
rect 1505 1937 1510 1942
rect 497 1932 550 1937
rect 577 1932 638 1937
rect 681 1932 742 1937
rect 753 1932 822 1937
rect 497 1927 502 1932
rect 481 1922 502 1927
rect 545 1927 550 1932
rect 545 1922 622 1927
rect 737 1922 742 1932
rect 817 1927 822 1932
rect 881 1932 926 1937
rect 1273 1932 1510 1937
rect 1697 1932 1822 1937
rect 881 1927 886 1932
rect 1953 1927 1958 1962
rect 817 1922 886 1927
rect 1169 1922 1254 1927
rect 1529 1922 1638 1927
rect 1649 1922 1814 1927
rect 1921 1922 1958 1927
rect 1169 1917 1174 1922
rect 497 1912 558 1917
rect 585 1912 614 1917
rect 657 1912 686 1917
rect 681 1907 686 1912
rect 761 1912 790 1917
rect 1145 1912 1174 1917
rect 1305 1912 1398 1917
rect 1561 1912 1598 1917
rect 1633 1912 1638 1922
rect 1689 1912 1910 1917
rect 761 1907 766 1912
rect 273 1902 374 1907
rect 681 1902 766 1907
rect 857 1902 998 1907
rect 1009 1902 1214 1907
rect 1841 1902 1910 1907
rect 257 1892 294 1897
rect 1889 1892 1974 1897
rect 1985 1887 1990 1957
rect 2153 1952 2230 1957
rect 2049 1942 2166 1947
rect 2345 1942 2510 1947
rect 2097 1932 2222 1937
rect 2073 1912 2126 1917
rect 2161 1912 2166 1932
rect 2225 1912 2278 1917
rect 2385 1912 2390 1937
rect 2409 1912 2598 1917
rect 2001 1902 2118 1907
rect 2137 1902 2254 1907
rect 2401 1902 2486 1907
rect 2017 1892 2070 1897
rect 2177 1892 2246 1897
rect 345 1882 366 1887
rect 433 1882 542 1887
rect 433 1867 438 1882
rect 537 1877 542 1882
rect 1329 1882 1478 1887
rect 1793 1882 1878 1887
rect 1985 1882 2014 1887
rect 2025 1882 2078 1887
rect 1329 1877 1334 1882
rect 537 1872 566 1877
rect 585 1872 750 1877
rect 1305 1872 1334 1877
rect 1473 1877 1478 1882
rect 1473 1872 1502 1877
rect 1849 1872 1878 1877
rect 241 1862 438 1867
rect 449 1862 478 1867
rect 585 1862 590 1872
rect 497 1857 590 1862
rect 745 1857 750 1872
rect 929 1862 1014 1867
rect 1329 1862 1486 1867
rect 2089 1862 2206 1867
rect 369 1852 502 1857
rect 745 1852 822 1857
rect 2105 1852 2214 1857
rect 177 1842 302 1847
rect 457 1842 518 1847
rect 537 1842 734 1847
rect 1425 1842 1542 1847
rect 2017 1842 2110 1847
rect 153 1832 286 1837
rect 297 1832 382 1837
rect 513 1827 518 1842
rect 1425 1837 1430 1842
rect 1369 1832 1430 1837
rect 1537 1837 1542 1842
rect 1537 1832 1566 1837
rect 1753 1832 1830 1837
rect 1857 1832 1926 1837
rect 2049 1832 2190 1837
rect 2369 1832 2422 1837
rect 2489 1832 2550 1837
rect 2593 1832 2622 1837
rect 1753 1827 1758 1832
rect 169 1822 318 1827
rect 513 1822 550 1827
rect 713 1822 782 1827
rect 977 1822 1022 1827
rect 1441 1822 1478 1827
rect 1489 1822 1574 1827
rect 1641 1822 1686 1827
rect 1729 1822 1758 1827
rect 1825 1827 1830 1832
rect 1825 1822 1854 1827
rect 1865 1822 1902 1827
rect 1937 1822 1982 1827
rect 2033 1822 2062 1827
rect 2169 1822 2214 1827
rect 2225 1822 2262 1827
rect 2337 1822 2406 1827
rect 2537 1822 2590 1827
rect 2601 1822 2646 1827
rect 137 1792 158 1797
rect 241 1782 246 1817
rect 257 1782 262 1817
rect 281 1812 310 1817
rect 337 1812 366 1817
rect 577 1812 670 1817
rect 761 1812 790 1817
rect 801 1812 838 1817
rect 1457 1812 1518 1817
rect 1777 1812 1894 1817
rect 1969 1812 2006 1817
rect 2073 1812 2198 1817
rect 2209 1807 2214 1822
rect 441 1802 494 1807
rect 521 1802 750 1807
rect 913 1802 998 1807
rect 1009 1802 1062 1807
rect 1705 1802 1798 1807
rect 2009 1802 2086 1807
rect 2169 1802 2214 1807
rect 297 1792 406 1797
rect 465 1792 606 1797
rect 1417 1792 1438 1797
rect 1465 1792 1510 1797
rect 1633 1792 1718 1797
rect 1745 1792 1790 1797
rect 2097 1792 2302 1797
rect 409 1782 526 1787
rect 601 1782 630 1787
rect 665 1782 710 1787
rect 921 1782 1086 1787
rect 1425 1782 1502 1787
rect 2017 1782 2062 1787
rect 2089 1782 2142 1787
rect 2177 1782 2262 1787
rect 2385 1777 2390 1817
rect 2425 1812 2606 1817
rect 2465 1802 2598 1807
rect 2425 1782 2502 1787
rect 2569 1782 2630 1787
rect 433 1772 686 1777
rect 817 1772 966 1777
rect 1313 1772 1398 1777
rect 1521 1772 1558 1777
rect 1713 1772 1790 1777
rect 2113 1772 2158 1777
rect 2345 1772 2390 1777
rect 2433 1772 2622 1777
rect 1313 1767 1318 1772
rect 441 1762 494 1767
rect 545 1762 654 1767
rect 1289 1762 1318 1767
rect 1393 1767 1398 1772
rect 1713 1767 1718 1772
rect 1785 1767 1862 1772
rect 1393 1762 1718 1767
rect 1857 1762 1998 1767
rect 2329 1762 2366 1767
rect 193 1752 222 1757
rect 377 1752 438 1757
rect 481 1752 582 1757
rect 593 1752 662 1757
rect 1033 1752 1118 1757
rect 1521 1752 1606 1757
rect 1729 1752 1774 1757
rect 105 1742 166 1747
rect 209 1742 326 1747
rect 441 1742 486 1747
rect 609 1742 646 1747
rect 993 1742 1070 1747
rect 1297 1742 1422 1747
rect 481 1737 486 1742
rect 465 1727 470 1737
rect 481 1732 622 1737
rect 681 1732 742 1737
rect 937 1732 1126 1737
rect 1233 1727 1238 1737
rect 1441 1732 1518 1737
rect 169 1722 222 1727
rect 409 1722 446 1727
rect 465 1722 486 1727
rect 497 1722 542 1727
rect 553 1722 622 1727
rect 633 1722 750 1727
rect 1049 1722 1158 1727
rect 1209 1722 1238 1727
rect 1313 1722 1382 1727
rect 1449 1722 1534 1727
rect 153 1712 182 1717
rect 441 1712 494 1717
rect 609 1712 670 1717
rect 857 1712 1046 1717
rect 1193 1712 1238 1717
rect 1409 1712 1446 1717
rect 1457 1712 1486 1717
rect 1641 1712 1678 1717
rect 1729 1707 1734 1752
rect 1841 1737 1846 1757
rect 2353 1752 2398 1757
rect 2433 1752 2494 1757
rect 2249 1742 2294 1747
rect 2377 1742 2574 1747
rect 1841 1732 1878 1737
rect 2129 1732 2222 1737
rect 2425 1732 2494 1737
rect 2529 1732 2566 1737
rect 1753 1722 1862 1727
rect 1873 1722 1878 1732
rect 2161 1722 2294 1727
rect 2449 1722 2486 1727
rect 1857 1717 1862 1722
rect 1761 1712 1798 1717
rect 1857 1712 1902 1717
rect 2145 1712 2206 1717
rect 2233 1712 2270 1717
rect 2473 1712 2502 1717
rect 121 1702 142 1707
rect 361 1702 438 1707
rect 465 1702 606 1707
rect 657 1702 766 1707
rect 1161 1702 1246 1707
rect 1329 1702 1358 1707
rect 1353 1697 1358 1702
rect 1433 1702 1494 1707
rect 1729 1702 1790 1707
rect 1809 1702 1846 1707
rect 2113 1702 2166 1707
rect 2201 1702 2262 1707
rect 2337 1702 2366 1707
rect 2425 1702 2510 1707
rect 2569 1702 2606 1707
rect 1433 1697 1438 1702
rect 561 1692 734 1697
rect 1353 1692 1438 1697
rect 1665 1692 1830 1697
rect 1841 1692 1878 1697
rect 2209 1692 2246 1697
rect 2465 1692 2638 1697
rect 1825 1687 1830 1692
rect 625 1682 710 1687
rect 1473 1682 1558 1687
rect 1585 1682 1782 1687
rect 1825 1682 1878 1687
rect 2321 1682 2358 1687
rect 2481 1682 2582 1687
rect 2601 1682 2646 1687
rect 1873 1677 1878 1682
rect 409 1672 542 1677
rect 753 1672 934 1677
rect 1457 1672 1550 1677
rect 1633 1672 1710 1677
rect 1873 1672 1966 1677
rect 2001 1672 2102 1677
rect 409 1667 414 1672
rect 537 1667 702 1672
rect 753 1667 758 1672
rect 185 1662 414 1667
rect 697 1662 758 1667
rect 929 1667 934 1672
rect 929 1662 958 1667
rect 1497 1662 1582 1667
rect 481 1652 686 1657
rect 825 1652 910 1657
rect 921 1652 942 1657
rect 1465 1652 1558 1657
rect 1729 1652 1854 1657
rect 1921 1652 1974 1657
rect 1985 1652 2006 1657
rect 705 1647 806 1652
rect 1729 1647 1734 1652
rect 209 1642 246 1647
rect 425 1642 526 1647
rect 601 1642 710 1647
rect 801 1642 998 1647
rect 1353 1642 1526 1647
rect 1593 1642 1654 1647
rect 1697 1642 1734 1647
rect 1849 1647 1854 1652
rect 1849 1642 2094 1647
rect 2513 1642 2550 1647
rect 993 1637 998 1642
rect 193 1632 286 1637
rect 297 1632 390 1637
rect 449 1632 558 1637
rect 641 1632 742 1637
rect 753 1632 934 1637
rect 993 1632 1110 1637
rect 1201 1632 1294 1637
rect 1409 1632 1510 1637
rect 1545 1632 1678 1637
rect 1745 1632 1814 1637
rect 1833 1632 1918 1637
rect 1745 1627 1750 1632
rect 1913 1627 1918 1632
rect 1985 1632 2014 1637
rect 2361 1632 2406 1637
rect 2465 1632 2526 1637
rect 1985 1627 1990 1632
rect 161 1622 254 1627
rect 281 1622 318 1627
rect 329 1622 358 1627
rect 377 1622 478 1627
rect 737 1622 782 1627
rect 889 1622 934 1627
rect 1025 1622 1126 1627
rect 321 1612 342 1617
rect 361 1612 406 1617
rect 521 1612 758 1617
rect 801 1612 854 1617
rect 865 1612 1174 1617
rect 265 1602 326 1607
rect 393 1602 494 1607
rect 721 1602 990 1607
rect 321 1597 326 1602
rect 1009 1597 1014 1612
rect 1185 1607 1190 1627
rect 1265 1622 1302 1627
rect 1313 1622 1422 1627
rect 1449 1622 1494 1627
rect 1521 1622 1622 1627
rect 1257 1612 1422 1617
rect 1433 1612 1558 1617
rect 1585 1612 1622 1617
rect 1169 1602 1190 1607
rect 1425 1602 1486 1607
rect 1169 1597 1174 1602
rect 1425 1597 1430 1602
rect 233 1592 310 1597
rect 321 1592 358 1597
rect 417 1592 542 1597
rect 569 1592 846 1597
rect 881 1592 982 1597
rect 1009 1592 1030 1597
rect 1105 1592 1174 1597
rect 1297 1592 1430 1597
rect 1489 1592 1566 1597
rect 1617 1587 1622 1612
rect 329 1582 358 1587
rect 393 1582 590 1587
rect 649 1582 694 1587
rect 705 1582 758 1587
rect 769 1582 838 1587
rect 993 1582 1190 1587
rect 1497 1582 1542 1587
rect 1593 1582 1622 1587
rect 1633 1582 1638 1617
rect 1649 1582 1654 1627
rect 1729 1622 1750 1627
rect 1761 1597 1766 1627
rect 1841 1622 1870 1627
rect 1913 1622 1990 1627
rect 2057 1622 2086 1627
rect 2105 1622 2142 1627
rect 2169 1622 2230 1627
rect 2257 1622 2318 1627
rect 2393 1622 2478 1627
rect 2497 1622 2590 1627
rect 1841 1617 1846 1622
rect 1777 1612 1846 1617
rect 1665 1592 1766 1597
rect 1673 1582 1726 1587
rect 1873 1582 1878 1617
rect 2081 1607 2086 1622
rect 2273 1612 2382 1617
rect 2401 1612 2454 1617
rect 2081 1602 2262 1607
rect 2345 1602 2374 1607
rect 2257 1597 2350 1602
rect 1913 1592 2022 1597
rect 1921 1582 1958 1587
rect 2153 1582 2198 1587
rect 2265 1582 2310 1587
rect 689 1577 694 1582
rect 769 1577 774 1582
rect 865 1577 998 1582
rect 1209 1577 1326 1582
rect 1385 1577 1478 1582
rect 345 1572 374 1577
rect 521 1572 606 1577
rect 689 1572 726 1577
rect 745 1572 774 1577
rect 809 1572 870 1577
rect 1017 1572 1046 1577
rect 1097 1572 1214 1577
rect 1321 1572 1390 1577
rect 1473 1572 1966 1577
rect 2281 1572 2438 1577
rect 369 1567 526 1572
rect 2497 1567 2502 1622
rect 2513 1612 2550 1617
rect 2577 1612 2598 1617
rect 2513 1582 2518 1612
rect 2537 1582 2566 1587
rect 2593 1582 2598 1612
rect 2609 1587 2614 1617
rect 2609 1582 2662 1587
rect 2545 1572 2606 1577
rect 545 1557 550 1567
rect 593 1562 718 1567
rect 737 1562 798 1567
rect 825 1562 926 1567
rect 953 1562 1110 1567
rect 1121 1562 1150 1567
rect 1177 1562 1214 1567
rect 1273 1562 1310 1567
rect 1401 1562 1526 1567
rect 1633 1562 1726 1567
rect 1929 1562 1958 1567
rect 2073 1562 2102 1567
rect 2233 1562 2334 1567
rect 2497 1562 2606 1567
rect 409 1552 462 1557
rect 481 1547 486 1557
rect 545 1552 558 1557
rect 577 1552 902 1557
rect 969 1552 1022 1557
rect 1057 1552 1102 1557
rect 1209 1552 1582 1557
rect 1601 1552 1678 1557
rect 1873 1552 1918 1557
rect 553 1547 558 1552
rect 1601 1547 1606 1552
rect 81 1542 182 1547
rect 361 1542 430 1547
rect 481 1542 542 1547
rect 553 1542 566 1547
rect 657 1542 710 1547
rect 361 1522 438 1527
rect 561 1522 566 1542
rect 737 1527 742 1547
rect 801 1527 806 1547
rect 961 1542 998 1547
rect 1201 1542 1262 1547
rect 1281 1542 1342 1547
rect 1377 1542 1406 1547
rect 1433 1542 1510 1547
rect 1561 1542 1606 1547
rect 1777 1542 1902 1547
rect 1377 1537 1382 1542
rect 897 1532 974 1537
rect 1321 1532 1382 1537
rect 1417 1532 1510 1537
rect 649 1522 790 1527
rect 801 1522 822 1527
rect 841 1522 1030 1527
rect 1113 1522 1174 1527
rect 1265 1522 1462 1527
rect 1505 1517 1510 1532
rect 1537 1517 1542 1527
rect 1657 1522 1686 1527
rect 1825 1522 1862 1527
rect 1953 1522 1958 1562
rect 1969 1547 1974 1557
rect 2025 1552 2142 1557
rect 2249 1552 2358 1557
rect 2481 1552 2534 1557
rect 2545 1547 2550 1557
rect 1969 1542 2070 1547
rect 2241 1542 2270 1547
rect 2265 1537 2270 1542
rect 2353 1542 2382 1547
rect 2497 1542 2550 1547
rect 2353 1537 2358 1542
rect 2089 1532 2214 1537
rect 2265 1532 2358 1537
rect 2441 1532 2526 1537
rect 2089 1527 2094 1532
rect 1993 1522 2094 1527
rect 2209 1527 2214 1532
rect 2609 1527 2614 1547
rect 2209 1522 2230 1527
rect 2385 1522 2430 1527
rect 2465 1522 2614 1527
rect 257 1512 310 1517
rect 545 1512 694 1517
rect 745 1512 838 1517
rect 857 1512 902 1517
rect 913 1512 942 1517
rect 1049 1512 1094 1517
rect 1289 1512 1326 1517
rect 1393 1512 1438 1517
rect 1481 1512 1510 1517
rect 1521 1512 1542 1517
rect 1713 1512 1750 1517
rect 1857 1512 1862 1522
rect 1961 1512 2054 1517
rect 2065 1512 2126 1517
rect 2145 1512 2206 1517
rect 2225 1512 2230 1522
rect 2409 1512 2438 1517
rect 2449 1512 2518 1517
rect 2553 1512 2646 1517
rect 161 1502 302 1507
rect 321 1502 414 1507
rect 601 1502 702 1507
rect 849 1502 1166 1507
rect 1425 1502 1542 1507
rect 1609 1502 1694 1507
rect 721 1497 830 1502
rect 1689 1497 1694 1502
rect 1761 1502 1806 1507
rect 1913 1502 1998 1507
rect 2081 1502 2358 1507
rect 2481 1502 2614 1507
rect 1761 1497 1766 1502
rect 681 1492 726 1497
rect 825 1492 982 1497
rect 1041 1492 1094 1497
rect 1313 1492 1670 1497
rect 1689 1492 1766 1497
rect 2129 1492 2166 1497
rect 2417 1492 2470 1497
rect 657 1482 854 1487
rect 945 1482 1070 1487
rect 1145 1482 1326 1487
rect 1905 1482 1998 1487
rect 2017 1482 2078 1487
rect 2505 1482 2550 1487
rect 1905 1477 1910 1482
rect 633 1472 710 1477
rect 1009 1472 1206 1477
rect 1881 1472 1910 1477
rect 1993 1477 1998 1482
rect 1993 1472 2030 1477
rect 1225 1462 1342 1467
rect 1769 1462 2054 1467
rect 2097 1462 2238 1467
rect 2257 1462 2358 1467
rect 1105 1457 1230 1462
rect 1337 1457 1342 1462
rect 2097 1457 2102 1462
rect 553 1452 758 1457
rect 865 1452 918 1457
rect 1081 1452 1110 1457
rect 1337 1452 1366 1457
rect 1473 1452 1622 1457
rect 1905 1452 1934 1457
rect 2025 1452 2102 1457
rect 2233 1457 2238 1462
rect 2233 1452 2278 1457
rect 1473 1447 1478 1452
rect 881 1442 942 1447
rect 1105 1442 1246 1447
rect 1305 1442 1374 1447
rect 1449 1442 1478 1447
rect 1617 1447 1622 1452
rect 1929 1447 2030 1452
rect 1617 1442 1646 1447
rect 2049 1442 2286 1447
rect 2305 1442 2374 1447
rect 2305 1437 2310 1442
rect 129 1432 158 1437
rect 745 1432 846 1437
rect 857 1432 926 1437
rect 977 1432 1150 1437
rect 1297 1432 1430 1437
rect 1577 1432 2134 1437
rect 2193 1432 2310 1437
rect 2369 1437 2374 1442
rect 2369 1432 2398 1437
rect 689 1422 758 1427
rect 825 1422 1054 1427
rect 145 1412 182 1417
rect 377 1412 398 1417
rect 153 1392 174 1397
rect 393 1392 454 1397
rect 529 1382 534 1417
rect 593 1412 734 1417
rect 777 1412 998 1417
rect 1033 1412 1062 1417
rect 1057 1397 1062 1412
rect 705 1392 854 1397
rect 929 1392 982 1397
rect 1057 1392 1086 1397
rect 1105 1387 1110 1427
rect 1121 1397 1126 1417
rect 1137 1407 1142 1427
rect 1161 1422 1190 1427
rect 1273 1422 1310 1427
rect 1329 1422 1494 1427
rect 1529 1422 1558 1427
rect 1593 1422 1630 1427
rect 2065 1422 2110 1427
rect 2257 1422 2278 1427
rect 2305 1422 2374 1427
rect 2473 1422 2518 1427
rect 2529 1422 2630 1427
rect 1137 1402 1158 1407
rect 1121 1392 1142 1397
rect 1033 1382 1110 1387
rect 913 1377 1014 1382
rect 433 1372 502 1377
rect 433 1367 438 1372
rect 409 1362 438 1367
rect 497 1367 502 1372
rect 553 1372 622 1377
rect 889 1372 918 1377
rect 1009 1372 1102 1377
rect 1153 1372 1158 1402
rect 1169 1382 1174 1417
rect 1185 1397 1190 1422
rect 1913 1417 2022 1422
rect 1201 1412 1350 1417
rect 1481 1412 1590 1417
rect 1889 1412 1918 1417
rect 2017 1412 2046 1417
rect 2169 1412 2222 1417
rect 1297 1402 1390 1407
rect 1433 1402 1470 1407
rect 1881 1402 1990 1407
rect 2057 1402 2166 1407
rect 1985 1397 2062 1402
rect 1185 1392 1206 1397
rect 1257 1392 1318 1397
rect 1457 1392 1566 1397
rect 2257 1387 2262 1422
rect 2273 1412 2302 1417
rect 2457 1412 2486 1417
rect 2273 1392 2278 1412
rect 2505 1402 2558 1407
rect 2449 1392 2526 1397
rect 1417 1382 1614 1387
rect 1985 1382 2038 1387
rect 2145 1382 2246 1387
rect 2257 1382 2294 1387
rect 1169 1372 1254 1377
rect 1481 1372 1502 1377
rect 1513 1372 1542 1377
rect 2025 1372 2246 1377
rect 553 1367 558 1372
rect 497 1362 558 1367
rect 617 1367 622 1372
rect 1345 1367 1462 1372
rect 617 1362 646 1367
rect 777 1362 822 1367
rect 833 1362 870 1367
rect 881 1362 1046 1367
rect 1169 1362 1246 1367
rect 1321 1362 1350 1367
rect 1457 1362 1726 1367
rect 2121 1362 2182 1367
rect 833 1357 838 1362
rect 2177 1357 2182 1362
rect 2273 1362 2302 1367
rect 2273 1357 2278 1362
rect 425 1352 486 1357
rect 785 1352 838 1357
rect 985 1352 1134 1357
rect 1177 1352 1214 1357
rect 1377 1352 1510 1357
rect 1777 1352 1854 1357
rect 1873 1352 1918 1357
rect 2017 1352 2046 1357
rect 2073 1352 2118 1357
rect 2129 1352 2158 1357
rect 2177 1352 2278 1357
rect 2385 1352 2518 1357
rect 513 1347 622 1352
rect 1777 1347 1782 1352
rect 129 1342 158 1347
rect 217 1342 414 1347
rect 497 1342 518 1347
rect 617 1342 702 1347
rect 873 1342 950 1347
rect 993 1342 1222 1347
rect 1369 1342 1446 1347
rect 1529 1342 1622 1347
rect 1753 1342 1782 1347
rect 1849 1347 1854 1352
rect 1849 1342 2118 1347
rect -1 1327 6 1328
rect -1 1322 0 1327
rect 5 1322 118 1327
rect 129 1322 134 1342
rect 409 1337 502 1342
rect 265 1332 318 1337
rect 521 1332 606 1337
rect 1033 1332 1222 1337
rect 1241 1332 1350 1337
rect 1409 1332 1598 1337
rect 1673 1332 1782 1337
rect 1865 1332 2014 1337
rect 1241 1327 1246 1332
rect 273 1322 318 1327
rect 361 1322 398 1327
rect 737 1322 1062 1327
rect 1185 1322 1246 1327
rect 1345 1327 1350 1332
rect 1345 1322 1662 1327
rect 1697 1322 1830 1327
rect 1889 1322 1910 1327
rect 1993 1322 2118 1327
rect 2129 1322 2134 1352
rect 2377 1342 2406 1347
rect 2425 1342 2502 1347
rect 2497 1332 2550 1337
rect 2497 1327 2502 1332
rect 2145 1322 2214 1327
rect 2481 1322 2502 1327
rect 2545 1322 2574 1327
rect 2593 1322 2598 1357
rect -1 1321 6 1322
rect 113 1317 118 1322
rect 1057 1317 1190 1322
rect 1697 1317 1702 1322
rect 2145 1317 2150 1322
rect 113 1312 222 1317
rect 473 1312 550 1317
rect 993 1312 1038 1317
rect 1209 1312 1342 1317
rect 1385 1312 1406 1317
rect 1481 1312 1574 1317
rect 1585 1312 1622 1317
rect 1665 1312 1702 1317
rect 1729 1312 1774 1317
rect 1817 1312 1894 1317
rect 1913 1312 1958 1317
rect 2025 1312 2070 1317
rect 2081 1312 2150 1317
rect 2193 1312 2238 1317
rect 2409 1312 2470 1317
rect 2497 1312 2582 1317
rect 2609 1312 2630 1317
rect 545 1307 550 1312
rect 817 1307 974 1312
rect 2609 1307 2614 1312
rect 177 1302 214 1307
rect 441 1302 470 1307
rect 497 1302 526 1307
rect 545 1302 574 1307
rect 793 1302 822 1307
rect 969 1302 1270 1307
rect 1409 1302 1438 1307
rect 1561 1302 1638 1307
rect 2041 1302 2070 1307
rect 2177 1302 2390 1307
rect 2457 1302 2486 1307
rect 2521 1302 2558 1307
rect 2569 1302 2614 1307
rect 1265 1297 1414 1302
rect 281 1292 302 1297
rect 801 1292 1086 1297
rect 1513 1292 1606 1297
rect 2513 1292 2598 1297
rect 1129 1287 1246 1292
rect 169 1282 286 1287
rect 801 1282 1134 1287
rect 1241 1282 1342 1287
rect 1337 1277 1342 1282
rect 1449 1282 1526 1287
rect 1545 1282 1614 1287
rect 1449 1277 1454 1282
rect -27 1274 -20 1275
rect -27 1269 -26 1274
rect -21 1273 6 1274
rect -21 1269 0 1273
rect -27 1268 -20 1269
rect -1 1268 0 1269
rect 5 1268 6 1273
rect 729 1272 830 1277
rect 993 1272 1070 1277
rect 1145 1272 1230 1277
rect 1337 1272 1454 1277
rect -1 1267 6 1268
rect 825 1267 998 1272
rect 489 1262 806 1267
rect 1017 1262 1166 1267
rect 1185 1262 1238 1267
rect 1521 1257 1526 1282
rect 1905 1272 2022 1277
rect 2145 1272 2182 1277
rect 2201 1272 2414 1277
rect 1625 1262 1822 1267
rect 2201 1262 2206 1272
rect 1625 1257 1630 1262
rect 2121 1257 2206 1262
rect 2409 1257 2414 1272
rect 769 1252 790 1257
rect 833 1252 950 1257
rect 977 1252 1030 1257
rect 1049 1252 1094 1257
rect 1185 1252 1318 1257
rect 1521 1252 1630 1257
rect 1737 1252 1766 1257
rect 1833 1252 2126 1257
rect 2409 1252 2542 1257
rect 1761 1247 1838 1252
rect 801 1242 846 1247
rect 873 1242 1262 1247
rect 2137 1242 2294 1247
rect 2393 1242 2414 1247
rect 169 1232 190 1237
rect 433 1232 454 1237
rect 465 1232 542 1237
rect 569 1232 654 1237
rect 841 1232 878 1237
rect 913 1232 1094 1237
rect 1289 1232 1350 1237
rect 1425 1232 1486 1237
rect 1777 1232 1806 1237
rect 1985 1232 2078 1237
rect 2393 1232 2446 1237
rect 113 1222 166 1227
rect 513 1222 558 1227
rect 753 1222 798 1227
rect 153 1212 190 1217
rect 561 1212 582 1217
rect 577 1202 582 1212
rect 689 1212 726 1217
rect 601 1202 630 1207
rect 129 1192 190 1197
rect 201 1192 270 1197
rect 321 1192 366 1197
rect 433 1192 478 1197
rect 561 1192 646 1197
rect 689 1187 694 1212
rect 737 1202 806 1207
rect 705 1192 822 1197
rect 321 1182 358 1187
rect 449 1182 510 1187
rect 617 1182 694 1187
rect 705 1182 742 1187
rect 761 1182 854 1187
rect 881 1182 886 1227
rect 905 1222 942 1227
rect 1025 1222 1086 1227
rect 1129 1222 1174 1227
rect 1241 1222 1286 1227
rect 1329 1222 1430 1227
rect 1457 1222 1566 1227
rect 1689 1222 1734 1227
rect 1809 1222 1838 1227
rect 1857 1222 1934 1227
rect 2089 1222 2126 1227
rect 2153 1222 2190 1227
rect 2353 1222 2390 1227
rect 2425 1222 2454 1227
rect 2497 1222 2526 1227
rect 945 1187 950 1217
rect 961 1202 1014 1207
rect 1025 1197 1030 1222
rect 1065 1212 1110 1217
rect 1009 1192 1030 1197
rect 945 1182 1046 1187
rect 1065 1182 1094 1187
rect 1105 1182 1110 1212
rect 1121 1212 1230 1217
rect 1577 1212 1966 1217
rect 2057 1212 2150 1217
rect 2273 1212 2366 1217
rect 1121 1202 1126 1212
rect 1225 1207 1582 1212
rect 1633 1202 1750 1207
rect 2025 1202 2158 1207
rect 2473 1202 2502 1207
rect 1769 1197 1862 1202
rect 2177 1197 2326 1202
rect 1217 1192 1350 1197
rect 1377 1192 1774 1197
rect 1857 1192 1886 1197
rect 1929 1192 2182 1197
rect 2321 1192 2350 1197
rect 2433 1192 2526 1197
rect 2545 1192 2566 1197
rect 1377 1182 1382 1192
rect 1737 1182 1814 1187
rect 1873 1182 1902 1187
rect 1961 1182 1998 1187
rect 2017 1182 2054 1187
rect 2137 1182 2334 1187
rect 1041 1177 1046 1182
rect 1401 1177 1718 1182
rect 2409 1177 2494 1182
rect 353 1172 430 1177
rect 529 1172 558 1177
rect 681 1172 910 1177
rect 953 1172 1022 1177
rect 1041 1172 1406 1177
rect 1713 1172 1758 1177
rect 1841 1172 1926 1177
rect 2009 1172 2414 1177
rect 2489 1172 2518 1177
rect 1753 1167 1846 1172
rect 1921 1167 1926 1172
rect 265 1162 382 1167
rect 457 1162 894 1167
rect 1009 1162 1038 1167
rect 1057 1162 1142 1167
rect 1345 1162 1734 1167
rect 1865 1162 1910 1167
rect 1921 1162 2086 1167
rect 2113 1162 2166 1167
rect 2257 1162 2286 1167
rect 2425 1162 2534 1167
rect 2161 1157 2262 1162
rect 49 1152 246 1157
rect 281 1152 318 1157
rect 369 1152 454 1157
rect 489 1152 638 1157
rect -13 1147 -6 1148
rect 49 1147 54 1152
rect -13 1142 -12 1147
rect -7 1142 54 1147
rect -13 1141 -6 1142
rect 241 1137 246 1152
rect 689 1147 694 1157
rect 337 1142 406 1147
rect 473 1142 502 1147
rect 585 1142 694 1147
rect 705 1152 774 1157
rect 785 1152 822 1157
rect 849 1152 1086 1157
rect 241 1132 422 1137
rect 441 1132 470 1137
rect 505 1132 542 1137
rect 569 1132 654 1137
rect 705 1127 710 1152
rect 745 1142 766 1147
rect 737 1132 790 1137
rect 65 1122 190 1127
rect 185 1117 190 1122
rect 257 1122 294 1127
rect 409 1122 446 1127
rect 489 1122 710 1127
rect 729 1122 758 1127
rect 785 1122 790 1132
rect 817 1122 822 1152
rect 1081 1147 1086 1152
rect 1233 1152 1382 1157
rect 1393 1152 1510 1157
rect 1609 1152 1638 1157
rect 1649 1152 1782 1157
rect 1793 1152 1838 1157
rect 1881 1152 1974 1157
rect 1233 1147 1238 1152
rect 881 1142 942 1147
rect 1081 1142 1238 1147
rect 1257 1142 1286 1147
rect 1433 1142 1718 1147
rect 1729 1142 1918 1147
rect 1281 1137 1438 1142
rect 1985 1137 1990 1157
rect 1457 1132 1814 1137
rect 1809 1127 1814 1132
rect 1921 1132 1990 1137
rect 2001 1137 2006 1157
rect 2001 1132 2022 1137
rect 961 1122 1062 1127
rect 1305 1122 1566 1127
rect 1665 1122 1798 1127
rect 1809 1122 1846 1127
rect 257 1117 262 1122
rect 185 1112 262 1117
rect 433 1112 462 1117
rect 497 1112 526 1117
rect 537 1112 574 1117
rect 633 1112 670 1117
rect 689 1112 742 1117
rect 833 1112 870 1117
rect 889 1112 918 1117
rect 1081 1112 1118 1117
rect 1489 1112 1550 1117
rect 1729 1112 1774 1117
rect 1793 1112 1798 1122
rect 1849 1112 1878 1117
rect 689 1107 694 1112
rect 281 1102 326 1107
rect 417 1102 694 1107
rect 745 1102 846 1107
rect 1073 1102 1310 1107
rect 1921 1102 1926 1132
rect 2017 1127 2022 1132
rect 1993 1122 2022 1127
rect 1961 1112 2022 1117
rect 2065 1107 2070 1157
rect 2081 1152 2126 1157
rect 2345 1152 2406 1157
rect 2481 1152 2574 1157
rect 2081 1122 2086 1152
rect 2153 1142 2174 1147
rect 2273 1142 2438 1147
rect 2473 1142 2526 1147
rect 2521 1137 2526 1142
rect 2585 1142 2630 1147
rect 2585 1137 2590 1142
rect 2097 1132 2126 1137
rect 2185 1132 2502 1137
rect 2521 1132 2590 1137
rect 2097 1122 2102 1132
rect 2121 1127 2190 1132
rect 2265 1122 2310 1127
rect 2393 1122 2438 1127
rect 2497 1122 2502 1132
rect 2185 1112 2230 1117
rect 2369 1112 2430 1117
rect 2481 1112 2582 1117
rect 2593 1112 2638 1117
rect 2481 1107 2486 1112
rect 2009 1102 2070 1107
rect 2345 1102 2486 1107
rect 2577 1107 2582 1112
rect 2577 1102 2606 1107
rect 2089 1097 2254 1102
rect 569 1092 734 1097
rect 809 1092 846 1097
rect 1385 1092 1734 1097
rect 1729 1087 1734 1092
rect 1817 1092 2094 1097
rect 2249 1092 2278 1097
rect 2409 1092 2478 1097
rect 2609 1092 2646 1097
rect 1817 1087 1822 1092
rect 161 1082 182 1087
rect 345 1082 374 1087
rect 1297 1082 1398 1087
rect 1673 1082 1710 1087
rect 1729 1082 1822 1087
rect 1913 1082 1942 1087
rect 2025 1082 2230 1087
rect 2289 1082 2454 1087
rect 2473 1082 2622 1087
rect 1937 1077 2030 1082
rect 2225 1077 2294 1082
rect 665 1072 750 1077
rect 1841 1072 1910 1077
rect 1905 1067 1910 1072
rect 2049 1072 2102 1077
rect 2161 1072 2206 1077
rect 2049 1067 2054 1072
rect 553 1062 654 1067
rect 729 1062 758 1067
rect 1273 1062 1326 1067
rect 1417 1062 1654 1067
rect 1905 1062 2054 1067
rect 2073 1062 2302 1067
rect 2369 1062 2398 1067
rect 649 1057 734 1062
rect 825 1052 926 1057
rect 825 1047 830 1052
rect 161 1042 294 1047
rect 577 1042 630 1047
rect 713 1042 790 1047
rect 801 1042 830 1047
rect 921 1047 926 1052
rect 1145 1052 1254 1057
rect 1313 1052 1342 1057
rect 1145 1047 1150 1052
rect 921 1042 950 1047
rect 1025 1042 1150 1047
rect 1249 1047 1254 1052
rect 1417 1047 1422 1062
rect 1649 1047 1654 1062
rect 1745 1052 1774 1057
rect 1817 1052 1886 1057
rect 2137 1052 2174 1057
rect 1249 1042 1422 1047
rect 1521 1042 1606 1047
rect 1649 1042 1734 1047
rect 1809 1042 2022 1047
rect 2129 1042 2246 1047
rect 1521 1037 1526 1042
rect 241 1032 278 1037
rect 433 1032 638 1037
rect 777 1032 878 1037
rect 897 1032 1070 1037
rect 1241 1032 1294 1037
rect 1305 1032 1358 1037
rect 1385 1032 1486 1037
rect 1497 1032 1526 1037
rect 1601 1037 1606 1042
rect 1729 1037 1814 1042
rect 1601 1032 1646 1037
rect 1833 1032 1902 1037
rect 1985 1032 2006 1037
rect 2033 1032 2086 1037
rect 2105 1032 2230 1037
rect 2561 1032 2598 1037
rect 129 1017 134 1027
rect 153 1022 190 1027
rect 297 1022 358 1027
rect 369 1022 406 1027
rect 73 1012 110 1017
rect 129 1012 238 1017
rect 281 1012 326 1017
rect 433 1012 454 1017
rect -1 1007 6 1008
rect 433 1007 438 1012
rect -1 1002 0 1007
rect 5 1002 70 1007
rect 169 1002 214 1007
rect 241 1002 318 1007
rect 433 1002 462 1007
rect -1 1001 6 1002
rect 65 997 70 1002
rect 497 997 502 1027
rect 585 1022 678 1027
rect 729 1022 870 1027
rect 977 1022 1006 1027
rect 1161 1022 1270 1027
rect 1297 1022 1534 1027
rect 977 1017 982 1022
rect 1585 1017 1590 1027
rect 1665 1022 1702 1027
rect 1785 1022 1830 1027
rect 1945 1022 1974 1027
rect 2057 1022 2094 1027
rect 2145 1022 2190 1027
rect 2201 1022 2270 1027
rect 2481 1022 2582 1027
rect 601 1012 646 1017
rect 649 1002 686 1007
rect 753 997 758 1017
rect 65 992 150 997
rect 201 992 318 997
rect 377 992 454 997
rect 473 992 502 997
rect 529 992 566 997
rect 617 992 726 997
rect 753 992 782 997
rect 73 982 110 987
rect 393 982 446 987
rect 465 982 526 987
rect 705 982 766 987
rect 801 982 806 1017
rect 817 977 822 1017
rect 889 1012 982 1017
rect 1057 1012 1254 1017
rect 1369 1012 1414 1017
rect 1121 1002 1150 1007
rect 1257 1002 1286 1007
rect 1297 1002 1318 1007
rect 865 997 1022 1002
rect 1145 997 1262 1002
rect 841 992 870 997
rect 1017 992 1046 997
rect 897 982 982 987
rect 193 972 254 977
rect 337 972 422 977
rect 529 972 574 977
rect 745 972 822 977
rect 977 977 982 982
rect 1057 982 1182 987
rect 1297 982 1302 1002
rect 1409 982 1414 1012
rect 1473 1007 1478 1017
rect 1505 1012 1542 1017
rect 1553 1012 1590 1017
rect 1609 1012 1638 1017
rect 1713 1012 1846 1017
rect 1881 1012 1918 1017
rect 2097 1012 2166 1017
rect 2281 1012 2390 1017
rect 2505 1012 2646 1017
rect 1473 1002 1526 1007
rect 1449 992 1510 997
rect 1521 987 1526 1002
rect 1481 982 1526 987
rect 1537 982 1542 1012
rect 1633 1007 1718 1012
rect 2161 1007 2286 1012
rect 2089 1002 2142 1007
rect 2361 1002 2382 1007
rect 2401 997 2518 1002
rect 1721 992 1838 997
rect 1937 992 2070 997
rect 1937 987 1942 992
rect 1617 982 1646 987
rect 1841 982 1942 987
rect 2065 987 2070 992
rect 2161 992 2262 997
rect 2353 992 2406 997
rect 2513 992 2542 997
rect 2161 987 2166 992
rect 2065 982 2166 987
rect 2257 987 2262 992
rect 2257 982 2510 987
rect 2561 982 2622 987
rect 1057 977 1062 982
rect 977 972 1062 977
rect 1225 972 1326 977
rect 1849 972 1894 977
rect 2001 972 2246 977
rect 2441 972 2558 977
rect 1649 967 1718 972
rect 2289 967 2422 972
rect 425 962 614 967
rect 825 962 958 967
rect 1241 962 1286 967
rect 1441 962 1654 967
rect 1713 962 1798 967
rect 1897 962 2158 967
rect 2169 962 2294 967
rect 2417 962 2606 967
rect 265 952 302 957
rect 321 952 406 957
rect 521 952 814 957
rect 1121 952 1206 957
rect 1273 952 1358 957
rect 1473 952 1502 957
rect 1665 952 1702 957
rect 2033 952 2078 957
rect 2113 952 2134 957
rect 1121 947 1126 952
rect 169 942 246 947
rect 369 942 414 947
rect 513 942 542 947
rect 681 942 806 947
rect 945 942 1014 947
rect 1097 942 1126 947
rect 1201 947 1206 952
rect 1201 942 1294 947
rect 1329 942 1374 947
rect 1641 942 1710 947
rect 1913 942 2070 947
rect 169 937 174 942
rect 145 932 174 937
rect 241 937 246 942
rect 2225 937 2230 957
rect 2305 952 2342 957
rect 2377 952 2430 957
rect 2249 942 2302 947
rect 2361 942 2390 947
rect 241 932 278 937
rect 545 932 670 937
rect 825 932 1054 937
rect 1073 932 1342 937
rect 1729 932 1894 937
rect 2225 932 2246 937
rect 665 927 750 932
rect 825 927 830 932
rect 1729 927 1734 932
rect 81 922 158 927
rect 553 922 574 927
rect 745 922 830 927
rect 1001 922 1142 927
rect 1193 922 1310 927
rect 1345 922 1398 927
rect 1425 922 1462 927
rect 1665 922 1734 927
rect 1889 927 1894 932
rect 1889 922 1934 927
rect 2041 922 2078 927
rect 2385 922 2390 942
rect 2593 927 2598 937
rect 2433 922 2502 927
rect 2593 922 2638 927
rect 1137 917 1142 922
rect 1457 917 1462 922
rect 121 912 174 917
rect 225 912 294 917
rect 577 912 630 917
rect 681 912 726 917
rect 993 912 1110 917
rect 1137 912 1246 917
rect 1393 912 1446 917
rect 1457 912 1510 917
rect 1529 912 1630 917
rect 1649 912 1734 917
rect 2185 912 2214 917
rect 2281 912 2398 917
rect 2513 912 2550 917
rect 1393 907 1398 912
rect 1529 907 1534 912
rect 601 902 702 907
rect 1001 902 1174 907
rect 1185 902 1230 907
rect 1241 902 1398 907
rect 1409 902 1534 907
rect 1625 907 1630 912
rect 1913 907 2006 912
rect 2065 907 2150 912
rect 1625 902 1918 907
rect 2001 902 2070 907
rect 2145 902 2174 907
rect 2329 902 2358 907
rect 2409 902 2470 907
rect 2529 902 2582 907
rect 361 892 438 897
rect 673 892 782 897
rect 1057 892 1086 897
rect 1081 887 1086 892
rect 1193 892 1222 897
rect 1233 892 1270 897
rect 1321 892 1430 897
rect 1481 892 1566 897
rect 1721 892 1782 897
rect 1929 892 1990 897
rect 1193 887 1198 892
rect 1985 887 1990 892
rect 2081 892 2278 897
rect 2081 887 2086 892
rect 2273 887 2278 892
rect 2409 892 2518 897
rect 2409 887 2414 892
rect 345 882 382 887
rect 1081 882 1198 887
rect 1385 882 1550 887
rect 1585 882 1702 887
rect 1697 877 1702 882
rect 1801 882 1910 887
rect 1985 882 2086 887
rect 2105 882 2150 887
rect 2193 882 2254 887
rect 2273 882 2414 887
rect 2497 882 2526 887
rect 1801 877 1806 882
rect 1449 872 1598 877
rect 1697 872 1806 877
rect 1905 877 1910 882
rect 1905 872 1958 877
rect 1313 867 1430 872
rect 873 862 958 867
rect 1289 862 1318 867
rect 1425 862 1646 867
rect 1745 862 1774 867
rect 1825 862 1966 867
rect 2433 862 2534 867
rect 873 857 878 862
rect 761 852 878 857
rect 953 857 958 862
rect 953 852 1038 857
rect 1137 852 1326 857
rect 1321 847 1326 852
rect 1385 852 1414 857
rect 1425 852 1822 857
rect 1385 847 1390 852
rect 209 842 302 847
rect 561 842 814 847
rect 1321 842 1390 847
rect 1529 842 1558 847
rect 1737 842 1878 847
rect 2241 842 2294 847
rect 209 837 214 842
rect 185 832 214 837
rect 297 837 302 842
rect 1553 837 1742 842
rect 297 832 326 837
rect 497 832 566 837
rect 665 832 710 837
rect 785 832 814 837
rect 889 832 942 837
rect 217 822 366 827
rect 385 822 422 827
rect 561 822 646 827
rect 689 822 726 827
rect 769 822 798 827
rect 921 822 1046 827
rect 1065 822 1142 827
rect 1169 822 1262 827
rect -1 817 6 818
rect -1 812 0 817
rect 5 812 174 817
rect -1 811 6 812
rect 281 802 350 807
rect 401 802 486 807
rect 625 802 726 807
rect 625 797 630 802
rect 129 792 190 797
rect 425 792 454 797
rect 609 792 630 797
rect 641 792 678 797
rect 601 782 686 787
rect 769 782 774 822
rect 817 812 1014 817
rect 897 802 990 807
rect 1009 792 1062 797
rect 1121 792 1174 797
rect 1297 782 1302 837
rect 1337 822 1478 827
rect 1505 822 1542 827
rect 1553 822 1598 827
rect 1657 822 1702 827
rect 1481 812 1566 817
rect 1617 812 1646 817
rect 1505 802 1614 807
rect 1745 797 1750 817
rect 1761 807 1766 837
rect 1817 832 1862 837
rect 2249 832 2278 837
rect 1777 822 1814 827
rect 2017 822 2070 827
rect 2121 822 2262 827
rect 2473 822 2598 827
rect 1801 812 1830 817
rect 1857 812 2006 817
rect 2097 812 2134 817
rect 2273 812 2366 817
rect 2577 812 2614 817
rect 1761 802 1798 807
rect 1345 792 1422 797
rect 1489 792 1542 797
rect 1721 792 1750 797
rect 1825 787 1830 812
rect 2089 802 2302 807
rect 1841 792 1870 797
rect 1913 792 1950 797
rect 2545 792 2614 797
rect 1313 782 1406 787
rect 1673 782 1718 787
rect 1737 782 1830 787
rect 1865 782 2118 787
rect 2129 782 2246 787
rect 2113 777 2118 782
rect 649 772 686 777
rect 793 772 830 777
rect 865 772 990 777
rect 1129 772 1182 777
rect 1225 772 1670 777
rect 1769 772 2102 777
rect 2113 772 2142 777
rect 2257 772 2398 777
rect 865 767 870 772
rect 217 762 302 767
rect 321 762 406 767
rect 833 762 870 767
rect 985 767 990 772
rect 2137 767 2262 772
rect 985 762 1070 767
rect 1249 762 1350 767
rect 1601 762 1686 767
rect 1849 762 1878 767
rect 1921 762 1998 767
rect 217 757 222 762
rect 193 752 222 757
rect 297 757 302 762
rect 297 752 326 757
rect 417 752 518 757
rect 897 752 918 757
rect 953 752 1142 757
rect 1169 752 1206 757
rect 1297 752 1366 757
rect 1513 752 1550 757
rect 2105 752 2150 757
rect 2161 752 2222 757
rect 2241 752 2326 757
rect 321 747 422 752
rect 2241 747 2246 752
rect 25 742 110 747
rect 129 742 190 747
rect 881 742 1062 747
rect 1193 742 1262 747
rect 1489 742 1518 747
rect 1537 742 1566 747
rect 1585 742 1670 747
rect 1729 742 2046 747
rect 2137 742 2174 747
rect 2217 742 2246 747
rect 2321 747 2326 752
rect 2481 752 2542 757
rect 2481 747 2486 752
rect 2321 742 2350 747
rect 2441 742 2486 747
rect 2601 742 2630 747
rect -1 737 6 738
rect 25 737 30 742
rect -1 732 0 737
rect 5 732 30 737
rect 105 737 110 742
rect 1345 737 1470 742
rect 1585 737 1590 742
rect 105 732 198 737
rect 209 732 278 737
rect 329 732 382 737
rect 489 732 510 737
rect 769 732 1182 737
rect -1 731 6 732
rect 1177 727 1182 732
rect 1249 732 1350 737
rect 1465 732 1590 737
rect 1665 737 1670 742
rect 1665 732 1694 737
rect 1777 732 1838 737
rect 2233 732 2278 737
rect 2337 732 2382 737
rect 2425 732 2598 737
rect 1249 727 1254 732
rect 481 722 502 727
rect 945 722 966 727
rect -1 717 6 718
rect -1 712 0 717
rect 5 712 54 717
rect 73 712 174 717
rect 865 712 918 717
rect 961 712 966 722
rect -1 711 6 712
rect 49 697 54 712
rect 1025 707 1030 727
rect 1177 722 1254 727
rect 1361 722 1678 727
rect 1105 712 1134 717
rect 1105 707 1110 712
rect 185 702 358 707
rect 377 702 478 707
rect 537 702 614 707
rect 841 702 862 707
rect 921 702 1110 707
rect 1129 707 1134 712
rect 1273 712 1318 717
rect 1369 712 1406 717
rect 1505 712 1558 717
rect 1273 707 1278 712
rect 1673 707 1678 722
rect 1841 722 1870 727
rect 2041 722 2142 727
rect 2193 722 2262 727
rect 2329 722 2366 727
rect 2385 722 2430 727
rect 2465 722 2502 727
rect 2625 722 2630 742
rect 1841 707 1846 722
rect 1905 712 1950 717
rect 2265 712 2326 717
rect 2337 712 2406 717
rect 2465 712 2470 722
rect 2585 712 2622 717
rect 1129 702 1278 707
rect 1297 702 1398 707
rect 1513 702 1550 707
rect 1561 702 1614 707
rect 1673 702 1846 707
rect 1993 702 2150 707
rect 2281 702 2414 707
rect 185 697 190 702
rect 49 692 190 697
rect 401 692 502 697
rect 809 692 838 697
rect 833 687 838 692
rect 913 692 942 697
rect 1033 692 1110 697
rect 2161 692 2214 697
rect 2313 692 2350 697
rect 2513 692 2590 697
rect 913 687 918 692
rect 465 682 486 687
rect 833 682 918 687
rect 1529 682 1654 687
rect 2081 682 2182 687
rect 521 672 758 677
rect -88 662 78 667
rect -88 643 -83 662
rect 521 657 526 672
rect 177 652 238 657
rect 313 652 470 657
rect 489 652 526 657
rect 753 657 758 672
rect 1537 662 1566 667
rect 1673 662 1726 667
rect 753 652 782 657
rect 801 652 926 657
rect -89 642 -82 643
rect -89 637 -88 642
rect -83 637 -82 642
rect 313 637 318 652
rect -89 636 -82 637
rect 289 632 318 637
rect 465 637 470 652
rect 801 647 806 652
rect 505 642 806 647
rect 921 647 926 652
rect 985 652 1134 657
rect 1473 652 1694 657
rect 2489 652 2574 657
rect 985 647 990 652
rect 921 642 990 647
rect 1129 647 1134 652
rect 2489 647 2494 652
rect 1129 642 1198 647
rect 1497 642 1654 647
rect 1825 642 1846 647
rect 2233 642 2286 647
rect 2465 642 2494 647
rect 2569 647 2574 652
rect 2569 642 2598 647
rect 465 632 494 637
rect 849 632 894 637
rect 1449 632 1630 637
rect 2121 632 2278 637
rect 2481 632 2526 637
rect 513 627 614 632
rect 273 622 334 627
rect 417 622 518 627
rect 609 622 638 627
rect 417 617 422 622
rect -88 612 86 617
rect 217 612 246 617
rect 345 612 422 617
rect 441 612 598 617
rect 737 612 758 617
rect -88 341 -83 612
rect 241 607 350 612
rect 129 602 206 607
rect 529 602 630 607
rect 673 602 710 607
rect 225 592 294 597
rect 353 592 398 597
rect 409 592 502 597
rect 529 587 534 602
rect 625 597 630 602
rect 569 592 614 597
rect 625 592 694 597
rect 737 592 742 612
rect 153 582 214 587
rect 209 577 214 582
rect 353 582 446 587
rect 481 582 534 587
rect 577 582 630 587
rect 657 582 806 587
rect 353 577 358 582
rect 817 577 822 627
rect 873 622 910 627
rect 1001 622 1038 627
rect 1065 622 1118 627
rect 1185 622 1286 627
rect 1305 622 1366 627
rect 1505 622 1598 627
rect 1873 622 1902 627
rect 1921 622 2022 627
rect 2225 622 2326 627
rect 2489 622 2638 627
rect 897 607 902 617
rect 1145 612 1230 617
rect 1425 612 1566 617
rect 1609 612 1638 617
rect 873 602 902 607
rect 1129 602 1190 607
rect 1465 602 1526 607
rect 1585 602 1606 607
rect 1649 602 1670 607
rect 841 592 870 597
rect 881 592 982 597
rect 1097 592 1190 597
rect 1225 592 1278 597
rect 1417 592 1446 597
rect 1657 592 1718 597
rect 1745 587 1750 617
rect 1769 612 1790 617
rect 1961 612 1990 617
rect 2193 612 2254 617
rect 2505 612 2582 617
rect 2337 602 2422 607
rect 2545 602 2606 607
rect 2337 597 2342 602
rect 1841 592 1934 597
rect 1993 592 2342 597
rect 2457 592 2534 597
rect 2545 592 2622 597
rect 833 582 862 587
rect 1665 582 1694 587
rect 1721 582 1750 587
rect 2393 582 2430 587
rect 2481 582 2526 587
rect 2577 582 2614 587
rect 81 572 190 577
rect 209 572 358 577
rect 457 572 774 577
rect 793 572 822 577
rect 849 572 1022 577
rect 1761 572 1790 577
rect 1825 572 1854 577
rect 1961 572 2038 577
rect 1961 567 1966 572
rect 401 562 430 567
rect 521 562 726 567
rect 777 562 878 567
rect 1009 562 1094 567
rect 1201 562 1342 567
rect 1785 562 1966 567
rect 2033 567 2038 572
rect 2089 572 2166 577
rect 2089 567 2094 572
rect 2033 562 2094 567
rect 2161 567 2166 572
rect 2161 562 2262 567
rect 577 552 790 557
rect 577 547 582 552
rect 961 547 966 557
rect 145 542 286 547
rect 481 542 582 547
rect 593 542 662 547
rect 689 542 830 547
rect 929 542 966 547
rect -1 537 6 538
rect -1 532 0 537
rect 5 532 70 537
rect 305 532 430 537
rect 449 532 646 537
rect 785 532 806 537
rect -1 531 6 532
rect 305 527 310 532
rect 281 522 310 527
rect 425 527 430 532
rect 425 522 710 527
rect 801 522 806 532
rect 929 522 934 542
rect 1009 517 1014 562
rect 1089 552 1366 557
rect 1409 552 1486 557
rect 1681 552 1710 557
rect 1681 547 1686 552
rect 1105 542 1142 547
rect 1209 542 1246 547
rect 1297 542 1358 547
rect 1377 542 1438 547
rect 1577 542 1686 547
rect 1697 542 1782 547
rect 1121 532 1158 537
rect 1185 532 1294 537
rect 1561 532 1590 537
rect 1185 527 1190 532
rect 1033 522 1102 527
rect 1145 522 1190 527
rect 1321 522 1358 527
rect 1441 522 1502 527
rect 1873 522 1878 557
rect 1897 552 1926 557
rect 1921 547 1926 552
rect 1985 552 2022 557
rect 2105 552 2150 557
rect 1985 547 1990 552
rect 2145 547 2150 552
rect 2249 552 2278 557
rect 2353 552 2382 557
rect 2249 547 2254 552
rect 1921 542 1990 547
rect 2009 542 2126 547
rect 2145 542 2254 547
rect 2289 542 2374 547
rect 2409 542 2510 547
rect 2097 522 2190 527
rect 2369 522 2502 527
rect 2537 522 2574 527
rect 2625 522 2646 527
rect 89 512 246 517
rect 321 512 350 517
rect 345 507 350 512
rect 457 512 486 517
rect 521 512 582 517
rect 721 512 862 517
rect 873 512 950 517
rect 1009 512 1030 517
rect 1153 512 1206 517
rect 1225 512 1294 517
rect 1465 512 1566 517
rect 1577 512 1686 517
rect 1769 512 1902 517
rect 2017 512 2102 517
rect 2137 512 2294 517
rect 2505 512 2550 517
rect 457 507 462 512
rect 345 502 462 507
rect 665 502 854 507
rect 865 502 910 507
rect 1025 502 1030 512
rect 2545 507 2550 512
rect 2625 507 2630 522
rect 1129 502 1246 507
rect 1425 502 1534 507
rect 1569 502 1670 507
rect 1897 502 1990 507
rect 2049 502 2094 507
rect 2497 502 2526 507
rect 2545 502 2630 507
rect 529 492 726 497
rect 721 487 726 492
rect 833 492 902 497
rect 929 492 1006 497
rect 1169 492 1302 497
rect 1489 492 1726 497
rect 2433 492 2478 497
rect 2489 492 2518 497
rect 833 487 838 492
rect 601 482 638 487
rect 673 482 702 487
rect 721 482 838 487
rect 921 482 1310 487
rect 1457 482 1718 487
rect 377 472 518 477
rect 889 472 1070 477
rect 1145 467 1310 472
rect 857 462 934 467
rect 1041 462 1150 467
rect 1305 462 1982 467
rect 1161 452 1294 457
rect 2433 452 2534 457
rect 2553 452 2630 457
rect 2433 447 2438 452
rect 369 442 558 447
rect 841 442 918 447
rect 977 442 1086 447
rect 1225 442 1278 447
rect 2265 442 2390 447
rect 2409 442 2438 447
rect 2529 447 2534 452
rect 2529 442 2574 447
rect 369 437 374 442
rect 345 432 374 437
rect 553 437 558 442
rect 2265 437 2270 442
rect 553 432 582 437
rect 897 432 998 437
rect 1185 432 1286 437
rect 1353 432 1454 437
rect 1473 432 1790 437
rect 1865 432 1966 437
rect 2017 432 2086 437
rect 2129 432 2214 437
rect 2241 432 2270 437
rect 2385 437 2390 442
rect 2385 432 2430 437
rect 2497 432 2566 437
rect 2585 432 2606 437
rect 65 422 174 427
rect 217 422 398 427
rect 305 412 550 417
rect 561 407 566 427
rect 737 422 846 427
rect 873 422 926 427
rect 977 422 1046 427
rect 1113 422 1238 427
rect 1505 417 1510 427
rect 1553 422 1606 427
rect 1761 417 1766 427
rect 1777 422 1854 427
rect 1849 417 1854 422
rect 1977 422 2110 427
rect 2121 422 2382 427
rect 2401 422 2478 427
rect 1977 417 1982 422
rect 825 412 862 417
rect 913 412 1006 417
rect 1161 412 1270 417
rect 1361 412 1390 417
rect 1505 412 1574 417
rect 1609 412 1662 417
rect 1761 412 1782 417
rect 329 402 366 407
rect 521 402 566 407
rect 673 402 710 407
rect 849 402 886 407
rect 961 402 1118 407
rect 1177 402 1206 407
rect 1369 402 1398 407
rect 1777 402 1782 412
rect 1809 397 1814 417
rect 1849 412 1982 417
rect 2001 412 2070 417
rect 2041 397 2110 402
rect 129 392 190 397
rect 217 392 238 397
rect 281 392 350 397
rect 513 392 1134 397
rect 1433 392 1574 397
rect 1649 392 1758 397
rect 1777 392 1814 397
rect 1833 392 2046 397
rect 2105 392 2134 397
rect 1649 387 1654 392
rect 337 382 382 387
rect 505 382 550 387
rect 561 382 670 387
rect 801 382 870 387
rect 985 382 1054 387
rect 1097 382 1174 387
rect 1345 382 1422 387
rect 1585 382 1654 387
rect 1753 387 1758 392
rect 2145 387 2150 417
rect 2177 412 2246 417
rect 2289 412 2326 417
rect 2465 412 2510 417
rect 2545 412 2566 417
rect 2305 402 2334 407
rect 2497 402 2654 407
rect 2305 397 2310 402
rect 2233 392 2310 397
rect 1753 382 1846 387
rect 1873 382 1902 387
rect 2057 382 2086 387
rect 2121 382 2150 387
rect 2289 382 2406 387
rect 1417 377 1590 382
rect 305 372 342 377
rect 553 372 918 377
rect 1025 372 1110 377
rect 1665 372 1774 377
rect 1809 372 2054 377
rect 913 367 982 372
rect 225 362 310 367
rect 529 362 574 367
rect 593 362 654 367
rect 761 362 902 367
rect 977 362 1062 367
rect 1377 362 1598 367
rect 1769 362 1878 367
rect 1889 362 1966 367
rect 2033 362 2070 367
rect 2345 362 2454 367
rect 649 357 766 362
rect 897 357 902 362
rect 281 352 438 357
rect 609 352 630 357
rect 785 352 886 357
rect 897 352 966 357
rect 1265 352 1310 357
rect 1617 352 1686 357
rect 2025 352 2062 357
rect 2377 352 2414 357
rect 2529 352 2598 357
rect 609 347 614 352
rect 1617 347 1622 352
rect 129 342 190 347
rect 321 342 350 347
rect -89 340 -82 341
rect -89 335 -88 340
rect -83 335 -82 340
rect -89 334 -82 335
rect -1 337 6 338
rect 345 337 350 342
rect 449 342 542 347
rect 577 342 614 347
rect 625 342 686 347
rect 841 342 894 347
rect 1113 342 1238 347
rect 1321 342 1438 347
rect 449 337 454 342
rect 1233 337 1326 342
rect 1433 337 1438 342
rect 1545 342 1622 347
rect 1681 347 1686 352
rect 1681 342 1830 347
rect 1849 342 1870 347
rect 2081 342 2134 347
rect 2241 342 2294 347
rect 2329 342 2374 347
rect 2385 342 2574 347
rect 1545 337 1550 342
rect -1 332 0 337
rect 5 332 182 337
rect 257 332 318 337
rect 345 332 454 337
rect 713 332 894 337
rect 913 332 1014 337
rect 1361 332 1414 337
rect 1433 332 1550 337
rect 1569 332 1606 337
rect 1625 332 1670 337
rect 1953 332 2094 337
rect 2313 332 2382 337
rect -1 331 6 332
rect 913 327 918 332
rect 729 322 758 327
rect 753 317 758 322
rect 833 322 918 327
rect 1009 327 1014 332
rect 1953 327 1958 332
rect 1009 322 1038 327
rect 1161 322 1198 327
rect 1257 322 1326 327
rect 1609 322 1694 327
rect 1713 322 1750 327
rect 1889 322 1958 327
rect 1969 322 2054 327
rect 2209 322 2486 327
rect 833 317 838 322
rect 753 312 838 317
rect 857 312 998 317
rect 1065 312 1094 317
rect 1137 312 1294 317
rect 1649 312 1710 317
rect 1857 312 2006 317
rect 2041 312 2070 317
rect 2081 312 2118 317
rect 2249 312 2318 317
rect 2329 312 2478 317
rect 993 307 1070 312
rect 217 302 430 307
rect 1201 302 1398 307
rect 1489 302 1590 307
rect 1921 302 2014 307
rect 2025 302 2102 307
rect 2217 302 2270 307
rect 2281 302 2334 307
rect 2425 302 2550 307
rect 1489 297 1494 302
rect 273 292 302 297
rect 297 287 302 292
rect 401 292 430 297
rect 961 292 1094 297
rect 401 287 406 292
rect 1089 287 1094 292
rect 1209 292 1238 297
rect 1385 292 1430 297
rect 1465 292 1494 297
rect 1585 297 1590 302
rect 1585 292 1662 297
rect 2017 292 2078 297
rect 2257 292 2302 297
rect 1209 287 1214 292
rect 297 282 406 287
rect 641 282 702 287
rect 1089 282 1214 287
rect 1681 282 1790 287
rect 2289 282 2350 287
rect 1313 277 1686 282
rect 1785 277 1790 282
rect 1241 272 1318 277
rect 1785 272 2142 277
rect 441 262 550 267
rect 561 262 1070 267
rect 1329 262 1774 267
rect 1057 252 1294 257
rect 1441 252 1630 257
rect 729 242 822 247
rect 1377 242 1718 247
rect 1793 242 1870 247
rect 1953 242 2174 247
rect 729 237 734 242
rect 425 232 734 237
rect 817 237 822 242
rect 1793 237 1798 242
rect 817 232 878 237
rect 961 232 1046 237
rect 1481 232 1574 237
rect 1625 232 1798 237
rect 1865 237 1870 242
rect 1865 232 1894 237
rect 1993 232 2046 237
rect 2193 232 2230 237
rect 2249 232 2278 237
rect 2409 232 2430 237
rect 745 222 862 227
rect 1065 222 1222 227
rect 1353 222 1414 227
rect 1473 222 1534 227
rect 1561 222 1598 227
rect 1617 222 1670 227
rect 1969 222 2022 227
rect 2097 222 2126 227
rect 2369 222 2406 227
rect 2097 217 2102 222
rect 2433 217 2438 227
rect 977 212 1006 217
rect 1193 212 1326 217
rect 1449 212 1494 217
rect 1529 212 1846 217
rect 1897 212 1982 217
rect 2025 212 2102 217
rect 2201 212 2286 217
rect 2321 212 2542 217
rect 897 202 1046 207
rect 1497 202 1782 207
rect 1849 202 1878 207
rect 1873 197 1878 202
rect 1953 202 1982 207
rect 2057 202 2086 207
rect 2209 202 2342 207
rect 2401 202 2614 207
rect 1953 197 1958 202
rect 2401 197 2406 202
rect 2609 197 2614 202
rect -80 192 70 197
rect 129 192 190 197
rect 305 192 334 197
rect 377 192 446 197
rect 505 192 566 197
rect 657 192 726 197
rect 809 192 894 197
rect 1009 192 1270 197
rect 1401 192 1526 197
rect 1585 192 1774 197
rect 1873 192 1958 197
rect 2073 192 2110 197
rect 2225 192 2310 197
rect 2321 192 2406 197
rect 2425 192 2462 197
rect 2481 192 2582 197
rect 2609 192 2630 197
rect -80 -157 -75 192
rect 449 182 550 187
rect 657 182 718 187
rect 993 182 1054 187
rect 1297 182 1382 187
rect 1601 182 1630 187
rect 1721 182 1750 187
rect 2089 182 2126 187
rect 2217 182 2334 187
rect 2441 182 2542 187
rect -1 177 6 178
rect 1297 177 1302 182
rect -1 172 0 177
rect 5 172 174 177
rect 281 172 390 177
rect 1273 172 1302 177
rect 1377 177 1382 182
rect 1377 172 1462 177
rect 2281 172 2342 177
rect -1 171 6 172
rect 281 167 286 172
rect 217 162 286 167
rect 385 167 390 172
rect 433 167 542 172
rect 2337 167 2342 172
rect 2409 172 2438 177
rect 2409 167 2414 172
rect 385 162 438 167
rect 537 162 566 167
rect 577 162 614 167
rect 761 162 878 167
rect 1025 162 1206 167
rect 1249 162 1350 167
rect 1417 162 1462 167
rect 1481 162 1702 167
rect 577 157 582 162
rect 1481 157 1486 162
rect 153 152 582 157
rect 593 152 750 157
rect 849 152 990 157
rect 105 142 158 147
rect 169 142 230 147
rect 321 142 382 147
rect 473 142 534 147
rect 561 142 598 147
rect 625 142 686 147
rect 729 142 766 147
rect 777 142 862 147
rect 705 132 734 137
rect 881 132 974 137
rect 729 127 886 132
rect 225 122 702 127
rect 473 112 510 117
rect 561 112 590 117
rect 585 97 590 112
rect 713 112 830 117
rect 945 112 998 117
rect 1057 112 1062 157
rect 1145 152 1486 157
rect 1697 157 1702 162
rect 1985 162 2070 167
rect 2273 162 2318 167
rect 2337 162 2414 167
rect 1985 157 1990 162
rect 1697 152 1990 157
rect 2065 157 2070 162
rect 2065 152 2182 157
rect 1137 142 1166 147
rect 1161 137 1166 142
rect 1233 142 1262 147
rect 1289 142 1366 147
rect 1377 142 1430 147
rect 1441 142 1686 147
rect 2001 142 2030 147
rect 1233 137 1238 142
rect 1441 137 1446 142
rect 1161 132 1238 137
rect 1321 132 1358 137
rect 1369 132 1446 137
rect 1465 132 1766 137
rect 2033 132 2110 137
rect 2249 132 2294 137
rect 1329 122 1390 127
rect 1441 122 1638 127
rect 1673 122 1726 127
rect 1769 122 1822 127
rect 1889 122 1926 127
rect 2201 122 2270 127
rect 1217 112 1302 117
rect 1345 112 1710 117
rect 713 97 718 112
rect 1217 107 1222 112
rect 977 102 1118 107
rect 1193 102 1222 107
rect 1297 107 1302 112
rect 1705 107 1710 112
rect 1833 112 1878 117
rect 1833 107 1838 112
rect 1297 102 1342 107
rect 1369 102 1398 107
rect 1393 97 1398 102
rect 1465 102 1494 107
rect 1545 102 1582 107
rect 1633 102 1686 107
rect 1705 102 1838 107
rect 1873 107 1878 112
rect 1937 112 2022 117
rect 1937 107 1942 112
rect 1873 102 1942 107
rect 2017 107 2022 112
rect 2089 112 2118 117
rect 2089 107 2094 112
rect 2017 102 2094 107
rect 1465 97 1470 102
rect 289 92 358 97
rect 585 92 718 97
rect 1033 92 1062 97
rect 1145 92 1174 97
rect 1201 92 1310 97
rect 1393 92 1470 97
rect 1057 87 1150 92
rect 1089 72 1118 77
rect 1113 67 1118 72
rect 1321 72 2294 77
rect 1321 67 1326 72
rect 1113 62 1326 67
rect 1034 -157 1041 -156
rect -80 -162 1035 -157
rect 1040 -162 1041 -157
rect 1034 -163 1041 -162
<< pad >>
rect -1 3654 41 3695
rect 285 3652 330 3692
rect 599 3654 645 3693
rect 914 3651 953 3687
rect 1202 3661 1243 3695
rect 1516 3658 1550 3691
rect 1804 3658 1846 3698
rect 2100 3642 2139 3681
rect 2404 3644 2450 3692
rect 2692 3641 2737 3686
rect -1017 2631 -982 2669
rect -1015 2337 -978 2372
rect 3727 2625 3753 2657
rect 3725 2342 3760 2374
rect -1020 2027 -989 2060
rect 3719 2030 3748 2063
rect -1015 1735 -982 1769
rect 3730 1742 3760 1770
rect -1018 1445 -986 1478
rect 3736 1432 3764 1459
rect -1030 1125 -1000 1157
rect 3723 1142 3756 1174
rect -1016 830 -989 854
rect 3728 849 3750 870
rect -1020 538 -996 563
rect 3731 545 3756 570
rect -1023 245 -998 269
rect 3726 240 3752 268
rect -1024 -67 -993 -38
rect 3728 -65 3756 -35
rect 14 -1069 40 -1044
rect 311 -1078 343 -1050
rect 609 -1079 639 -1052
rect 914 -1072 941 -1046
rect 1205 -1055 1224 -1038
rect 1511 -1076 1536 -1053
rect 1816 -1074 1846 -1048
rect 2110 -1091 2138 -1067
rect 2418 -1094 2446 -1066
rect 2713 -1085 2736 -1061
use top_mod_new_VIA1  top_mod_new_VIA1_0
timestamp 1681708930
transform 1 0 24 0 1 2617
box -10 -10 10 10
use top_mod_new_VIA1  top_mod_new_VIA1_1
timestamp 1681708930
transform 1 0 2712 0 1 2617
box -10 -10 10 10
use top_mod_new_VIA1  top_mod_new_VIA1_2
timestamp 1681708930
transform 1 0 48 0 1 2593
box -10 -10 10 10
use M3_M2  M3_M2_0
timestamp 1681708930
transform 1 0 1332 0 1 2585
box -3 -3 3 3
use top_mod_new_VIA1  top_mod_new_VIA1_3
timestamp 1681708930
transform 1 0 2688 0 1 2593
box -10 -10 10 10
use top_mod_new_VIA0  top_mod_new_VIA0_0
timestamp 1681708930
transform 1 0 48 0 1 2570
box -10 -3 10 3
use M3_M2  M3_M2_20
timestamp 1681708930
transform 1 0 180 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4
timestamp 1681708930
transform 1 0 180 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_21
timestamp 1681708930
transform 1 0 276 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_5
timestamp 1681708930
transform 1 0 276 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_22
timestamp 1681708930
transform 1 0 372 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1
timestamp 1681708930
transform 1 0 564 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_23
timestamp 1681708930
transform 1 0 484 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_6
timestamp 1681708930
transform 1 0 372 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_44
timestamp 1681708930
transform 1 0 452 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_7
timestamp 1681708930
transform 1 0 460 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_8
timestamp 1681708930
transform 1 0 484 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_9
timestamp 1681708930
transform 1 0 580 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_24
timestamp 1681708930
transform 1 0 628 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_9
timestamp 1681708930
transform 1 0 580 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_25
timestamp 1681708930
transform 1 0 684 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_10
timestamp 1681708930
transform 1 0 684 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_70
timestamp 1681708930
transform 1 0 228 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_71
timestamp 1681708930
transform 1 0 260 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_72
timestamp 1681708930
transform 1 0 316 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_73
timestamp 1681708930
transform 1 0 356 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_74
timestamp 1681708930
transform 1 0 396 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_75
timestamp 1681708930
transform 1 0 452 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_76
timestamp 1681708930
transform 1 0 468 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_77
timestamp 1681708930
transform 1 0 508 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_78
timestamp 1681708930
transform 1 0 564 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_79
timestamp 1681708930
transform 1 0 628 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_80
timestamp 1681708930
transform 1 0 668 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_69
timestamp 1681708930
transform 1 0 228 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_70
timestamp 1681708930
transform 1 0 276 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_107
timestamp 1681708930
transform 1 0 356 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_91
timestamp 1681708930
transform 1 0 476 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_108
timestamp 1681708930
transform 1 0 556 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_71
timestamp 1681708930
transform 1 0 668 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_127
timestamp 1681708930
transform 1 0 684 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_92
timestamp 1681708930
transform 1 0 684 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_26
timestamp 1681708930
transform 1 0 716 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_11
timestamp 1681708930
transform 1 0 716 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_81
timestamp 1681708930
transform 1 0 724 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_12
timestamp 1681708930
transform 1 0 732 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_53
timestamp 1681708930
transform 1 0 732 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_13
timestamp 1681708930
transform 1 0 756 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_14
timestamp 1681708930
transform 1 0 772 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_82
timestamp 1681708930
transform 1 0 748 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_83
timestamp 1681708930
transform 1 0 764 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_128
timestamp 1681708930
transform 1 0 732 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_83
timestamp 1681708930
transform 1 0 724 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_84
timestamp 1681708930
transform 1 0 764 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2
timestamp 1681708930
transform 1 0 820 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_10
timestamp 1681708930
transform 1 0 804 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_27
timestamp 1681708930
transform 1 0 820 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_15
timestamp 1681708930
transform 1 0 804 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_16
timestamp 1681708930
transform 1 0 820 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4
timestamp 1681708930
transform 1 0 860 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5
timestamp 1681708930
transform 1 0 924 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_11
timestamp 1681708930
transform 1 0 852 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_28
timestamp 1681708930
transform 1 0 844 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_29
timestamp 1681708930
transform 1 0 884 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_17
timestamp 1681708930
transform 1 0 844 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_18
timestamp 1681708930
transform 1 0 860 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_19
timestamp 1681708930
transform 1 0 948 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_84
timestamp 1681708930
transform 1 0 828 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_54
timestamp 1681708930
transform 1 0 860 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_85
timestamp 1681708930
transform 1 0 884 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_86
timestamp 1681708930
transform 1 0 940 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_129
timestamp 1681708930
transform 1 0 844 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_93
timestamp 1681708930
transform 1 0 884 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_20
timestamp 1681708930
transform 1 0 964 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_87
timestamp 1681708930
transform 1 0 956 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3
timestamp 1681708930
transform 1 0 1092 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_6
timestamp 1681708930
transform 1 0 988 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_7
timestamp 1681708930
transform 1 0 1044 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1681708930
transform 1 0 1076 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_30
timestamp 1681708930
transform 1 0 1036 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_12
timestamp 1681708930
transform 1 0 1092 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_21
timestamp 1681708930
transform 1 0 988 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_22
timestamp 1681708930
transform 1 0 1076 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_23
timestamp 1681708930
transform 1 0 1092 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_88
timestamp 1681708930
transform 1 0 972 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_89
timestamp 1681708930
transform 1 0 1036 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_90
timestamp 1681708930
transform 1 0 1076 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_94
timestamp 1681708930
transform 1 0 1060 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_55
timestamp 1681708930
transform 1 0 1084 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_31
timestamp 1681708930
transform 1 0 1116 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_24
timestamp 1681708930
transform 1 0 1116 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_25
timestamp 1681708930
transform 1 0 1124 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_26
timestamp 1681708930
transform 1 0 1148 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_91
timestamp 1681708930
transform 1 0 1100 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_56
timestamp 1681708930
transform 1 0 1124 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_130
timestamp 1681708930
transform 1 0 1140 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_95
timestamp 1681708930
transform 1 0 1140 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_13
timestamp 1681708930
transform 1 0 1164 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_27
timestamp 1681708930
transform 1 0 1164 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_32
timestamp 1681708930
transform 1 0 1196 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_28
timestamp 1681708930
transform 1 0 1196 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_92
timestamp 1681708930
transform 1 0 1172 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_93
timestamp 1681708930
transform 1 0 1180 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_94
timestamp 1681708930
transform 1 0 1196 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_131
timestamp 1681708930
transform 1 0 1196 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_14
timestamp 1681708930
transform 1 0 1324 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_15
timestamp 1681708930
transform 1 0 1348 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_16
timestamp 1681708930
transform 1 0 1380 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_33
timestamp 1681708930
transform 1 0 1252 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_34
timestamp 1681708930
transform 1 0 1308 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_29
timestamp 1681708930
transform 1 0 1212 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_30
timestamp 1681708930
transform 1 0 1228 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_96
timestamp 1681708930
transform 1 0 1204 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_31
timestamp 1681708930
transform 1 0 1324 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_32
timestamp 1681708930
transform 1 0 1332 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_33
timestamp 1681708930
transform 1 0 1380 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_34
timestamp 1681708930
transform 1 0 1388 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_95
timestamp 1681708930
transform 1 0 1252 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_96
timestamp 1681708930
transform 1 0 1308 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_97
timestamp 1681708930
transform 1 0 1332 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_98
timestamp 1681708930
transform 1 0 1356 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_17
timestamp 1681708930
transform 1 0 1444 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_35
timestamp 1681708930
transform 1 0 1436 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_35
timestamp 1681708930
transform 1 0 1436 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_36
timestamp 1681708930
transform 1 0 1444 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1681708930
transform 1 0 1412 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_72
timestamp 1681708930
transform 1 0 1380 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_73
timestamp 1681708930
transform 1 0 1412 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_85
timestamp 1681708930
transform 1 0 1356 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_109
timestamp 1681708930
transform 1 0 1388 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_36
timestamp 1681708930
transform 1 0 1492 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_37
timestamp 1681708930
transform 1 0 1492 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_100
timestamp 1681708930
transform 1 0 1468 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_38
timestamp 1681708930
transform 1 0 1548 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_39
timestamp 1681708930
transform 1 0 1556 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_101
timestamp 1681708930
transform 1 0 1532 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_40
timestamp 1681708930
transform 1 0 1604 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_102
timestamp 1681708930
transform 1 0 1580 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_57
timestamp 1681708930
transform 1 0 1604 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_41
timestamp 1681708930
transform 1 0 1660 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_103
timestamp 1681708930
transform 1 0 1636 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_97
timestamp 1681708930
transform 1 0 1580 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_74
timestamp 1681708930
transform 1 0 1636 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_37
timestamp 1681708930
transform 1 0 1716 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_42
timestamp 1681708930
transform 1 0 1716 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_43
timestamp 1681708930
transform 1 0 1724 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1681708930
transform 1 0 1692 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_105
timestamp 1681708930
transform 1 0 1700 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_98
timestamp 1681708930
transform 1 0 1700 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_110
timestamp 1681708930
transform 1 0 1692 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_58
timestamp 1681708930
transform 1 0 1724 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_75
timestamp 1681708930
transform 1 0 1724 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_0
timestamp 1681708930
transform 1 0 1828 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_44
timestamp 1681708930
transform 1 0 1780 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_45
timestamp 1681708930
transform 1 0 1804 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_46
timestamp 1681708930
transform 1 0 1812 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_45
timestamp 1681708930
transform 1 0 1828 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_106
timestamp 1681708930
transform 1 0 1772 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_107
timestamp 1681708930
transform 1 0 1788 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_108
timestamp 1681708930
transform 1 0 1812 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_76
timestamp 1681708930
transform 1 0 1780 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_99
timestamp 1681708930
transform 1 0 1772 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_100
timestamp 1681708930
transform 1 0 1796 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_38
timestamp 1681708930
transform 1 0 1852 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_47
timestamp 1681708930
transform 1 0 1852 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_109
timestamp 1681708930
transform 1 0 1844 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_101
timestamp 1681708930
transform 1 0 1844 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_48
timestamp 1681708930
transform 1 0 1892 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_110
timestamp 1681708930
transform 1 0 1868 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_59
timestamp 1681708930
transform 1 0 1884 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_111
timestamp 1681708930
transform 1 0 1892 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_132
timestamp 1681708930
transform 1 0 1860 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_77
timestamp 1681708930
transform 1 0 1868 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_133
timestamp 1681708930
transform 1 0 1884 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_102
timestamp 1681708930
transform 1 0 1876 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_1
timestamp 1681708930
transform 1 0 1908 0 1 2545
box -2 -2 2 2
use M3_M2  M3_M2_46
timestamp 1681708930
transform 1 0 1908 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_47
timestamp 1681708930
transform 1 0 1924 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_49
timestamp 1681708930
transform 1 0 1948 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_112
timestamp 1681708930
transform 1 0 1932 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_103
timestamp 1681708930
transform 1 0 1932 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_113
timestamp 1681708930
transform 1 0 1972 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_60
timestamp 1681708930
transform 1 0 1980 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_134
timestamp 1681708930
transform 1 0 1980 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_50
timestamp 1681708930
transform 1 0 2012 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_51
timestamp 1681708930
transform 1 0 2020 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_48
timestamp 1681708930
transform 1 0 2028 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_52
timestamp 1681708930
transform 1 0 2036 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_114
timestamp 1681708930
transform 1 0 2036 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_135
timestamp 1681708930
transform 1 0 2036 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_39
timestamp 1681708930
transform 1 0 2100 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_53
timestamp 1681708930
transform 1 0 2092 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_54
timestamp 1681708930
transform 1 0 2100 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_55
timestamp 1681708930
transform 1 0 2164 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_56
timestamp 1681708930
transform 1 0 2172 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1681708930
transform 1 0 2132 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_116
timestamp 1681708930
transform 1 0 2180 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_104
timestamp 1681708930
transform 1 0 2172 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_111
timestamp 1681708930
transform 1 0 2172 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_40
timestamp 1681708930
transform 1 0 2252 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_57
timestamp 1681708930
transform 1 0 2252 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_49
timestamp 1681708930
transform 1 0 2284 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_41
timestamp 1681708930
transform 1 0 2316 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_58
timestamp 1681708930
transform 1 0 2292 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_59
timestamp 1681708930
transform 1 0 2300 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_50
timestamp 1681708930
transform 1 0 2308 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_60
timestamp 1681708930
transform 1 0 2316 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_117
timestamp 1681708930
transform 1 0 2276 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_118
timestamp 1681708930
transform 1 0 2292 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_86
timestamp 1681708930
transform 1 0 2268 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_61
timestamp 1681708930
transform 1 0 2300 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_51
timestamp 1681708930
transform 1 0 2348 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_119
timestamp 1681708930
transform 1 0 2332 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_136
timestamp 1681708930
transform 1 0 2300 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_137
timestamp 1681708930
transform 1 0 2324 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_42
timestamp 1681708930
transform 1 0 2380 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_61
timestamp 1681708930
transform 1 0 2380 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1681708930
transform 1 0 2356 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_62
timestamp 1681708930
transform 1 0 2372 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_138
timestamp 1681708930
transform 1 0 2340 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1681708930
transform 1 0 2348 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_78
timestamp 1681708930
transform 1 0 2364 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_140
timestamp 1681708930
transform 1 0 2372 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_87
timestamp 1681708930
transform 1 0 2340 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_144
timestamp 1681708930
transform 1 0 2364 0 1 2505
box -2 -2 2 2
use M3_M2  M3_M2_105
timestamp 1681708930
transform 1 0 2356 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_18
timestamp 1681708930
transform 1 0 2404 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_2
timestamp 1681708930
transform 1 0 2404 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_62
timestamp 1681708930
transform 1 0 2412 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1681708930
transform 1 0 2404 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_19
timestamp 1681708930
transform 1 0 2452 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_63
timestamp 1681708930
transform 1 0 2436 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_64
timestamp 1681708930
transform 1 0 2452 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_65
timestamp 1681708930
transform 1 0 2468 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1681708930
transform 1 0 2420 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_63
timestamp 1681708930
transform 1 0 2428 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_43
timestamp 1681708930
transform 1 0 2500 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_66
timestamp 1681708930
transform 1 0 2492 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_123
timestamp 1681708930
transform 1 0 2444 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_64
timestamp 1681708930
transform 1 0 2468 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_124
timestamp 1681708930
transform 1 0 2476 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_65
timestamp 1681708930
transform 1 0 2484 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_79
timestamp 1681708930
transform 1 0 2412 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_80
timestamp 1681708930
transform 1 0 2428 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_81
timestamp 1681708930
transform 1 0 2444 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_88
timestamp 1681708930
transform 1 0 2420 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_106
timestamp 1681708930
transform 1 0 2436 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_141
timestamp 1681708930
transform 1 0 2484 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_89
timestamp 1681708930
transform 1 0 2476 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_3
timestamp 1681708930
transform 1 0 2532 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_67
timestamp 1681708930
transform 1 0 2524 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_68
timestamp 1681708930
transform 1 0 2540 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_66
timestamp 1681708930
transform 1 0 2508 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_125
timestamp 1681708930
transform 1 0 2516 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_142
timestamp 1681708930
transform 1 0 2508 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_145
timestamp 1681708930
transform 1 0 2500 0 1 2505
box -2 -2 2 2
use M3_M2  M3_M2_90
timestamp 1681708930
transform 1 0 2508 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_52
timestamp 1681708930
transform 1 0 2548 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_67
timestamp 1681708930
transform 1 0 2532 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_126
timestamp 1681708930
transform 1 0 2540 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_82
timestamp 1681708930
transform 1 0 2540 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_68
timestamp 1681708930
transform 1 0 2564 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_143
timestamp 1681708930
transform 1 0 2564 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_69
timestamp 1681708930
transform 1 0 2628 0 1 2535
box -2 -2 2 2
use top_mod_new_VIA0  top_mod_new_VIA0_1
timestamp 1681708930
transform 1 0 2688 0 1 2570
box -10 -3 10 3
use top_mod_new_VIA0  top_mod_new_VIA0_2
timestamp 1681708930
transform 1 0 24 0 1 2470
box -10 -3 10 3
use FILL  FILL_0
timestamp 1681708930
transform 1 0 72 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1
timestamp 1681708930
transform 1 0 80 0 -1 2570
box -8 -3 16 105
use FILL  FILL_2
timestamp 1681708930
transform 1 0 88 0 -1 2570
box -8 -3 16 105
use FILL  FILL_3
timestamp 1681708930
transform 1 0 96 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4
timestamp 1681708930
transform 1 0 104 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5
timestamp 1681708930
transform 1 0 112 0 -1 2570
box -8 -3 16 105
use FILL  FILL_6
timestamp 1681708930
transform 1 0 120 0 -1 2570
box -8 -3 16 105
use FILL  FILL_7
timestamp 1681708930
transform 1 0 128 0 -1 2570
box -8 -3 16 105
use FILL  FILL_8
timestamp 1681708930
transform 1 0 136 0 -1 2570
box -8 -3 16 105
use FILL  FILL_9
timestamp 1681708930
transform 1 0 144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_10
timestamp 1681708930
transform 1 0 152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_11
timestamp 1681708930
transform 1 0 160 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_0
timestamp 1681708930
transform 1 0 168 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_1
timestamp 1681708930
transform 1 0 264 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_2
timestamp 1681708930
transform 1 0 360 0 -1 2570
box -8 -3 104 105
use M3_M2  M3_M2_112
timestamp 1681708930
transform 1 0 468 0 1 2475
box -3 -3 3 3
use INVX2  INVX2_0
timestamp 1681708930
transform 1 0 456 0 -1 2570
box -9 -3 26 105
use M3_M2  M3_M2_113
timestamp 1681708930
transform 1 0 492 0 1 2475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_3
timestamp 1681708930
transform 1 0 472 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_4
timestamp 1681708930
transform 1 0 568 0 -1 2570
box -8 -3 104 105
use NAND2X1  NAND2X1_0
timestamp 1681708930
transform 1 0 664 0 -1 2570
box -8 -3 32 105
use OAI21X1  OAI21X1_0
timestamp 1681708930
transform -1 0 720 0 -1 2570
box -8 -3 34 105
use FILL  FILL_12
timestamp 1681708930
transform 1 0 720 0 -1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_1
timestamp 1681708930
transform -1 0 760 0 -1 2570
box -8 -3 34 105
use INVX2  INVX2_1
timestamp 1681708930
transform -1 0 776 0 -1 2570
box -9 -3 26 105
use FILL  FILL_13
timestamp 1681708930
transform 1 0 776 0 -1 2570
box -8 -3 16 105
use FILL  FILL_14
timestamp 1681708930
transform 1 0 784 0 -1 2570
box -8 -3 16 105
use FILL  FILL_15
timestamp 1681708930
transform 1 0 792 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_2
timestamp 1681708930
transform 1 0 800 0 -1 2570
box -9 -3 26 105
use OAI21X1  OAI21X1_2
timestamp 1681708930
transform 1 0 816 0 -1 2570
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_5
timestamp 1681708930
transform 1 0 848 0 -1 2570
box -8 -3 104 105
use INVX2  INVX2_3
timestamp 1681708930
transform 1 0 944 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_4
timestamp 1681708930
transform 1 0 960 0 -1 2570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_6
timestamp 1681708930
transform 1 0 976 0 -1 2570
box -8 -3 104 105
use INVX2  INVX2_5
timestamp 1681708930
transform 1 0 1072 0 -1 2570
box -9 -3 26 105
use OAI21X1  OAI21X1_3
timestamp 1681708930
transform 1 0 1088 0 -1 2570
box -8 -3 34 105
use M3_M2  M3_M2_114
timestamp 1681708930
transform 1 0 1148 0 1 2475
box -3 -3 3 3
use NAND2X1  NAND2X1_1
timestamp 1681708930
transform 1 0 1120 0 -1 2570
box -8 -3 32 105
use INVX2  INVX2_6
timestamp 1681708930
transform 1 0 1144 0 -1 2570
box -9 -3 26 105
use FILL  FILL_16
timestamp 1681708930
transform 1 0 1160 0 -1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_4
timestamp 1681708930
transform 1 0 1168 0 -1 2570
box -8 -3 34 105
use INVX2  INVX2_7
timestamp 1681708930
transform -1 0 1216 0 -1 2570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_7
timestamp 1681708930
transform 1 0 1216 0 -1 2570
box -8 -3 104 105
use INVX2  INVX2_8
timestamp 1681708930
transform -1 0 1328 0 -1 2570
box -9 -3 26 105
use XOR2X1  XOR2X1_0
timestamp 1681708930
transform -1 0 1384 0 -1 2570
box -8 -3 64 105
use XOR2X1  XOR2X1_1
timestamp 1681708930
transform -1 0 1440 0 -1 2570
box -8 -3 64 105
use XOR2X1  XOR2X1_2
timestamp 1681708930
transform -1 0 1496 0 -1 2570
box -8 -3 64 105
use M3_M2  M3_M2_115
timestamp 1681708930
transform 1 0 1556 0 1 2475
box -3 -3 3 3
use XOR2X1  XOR2X1_3
timestamp 1681708930
transform 1 0 1496 0 -1 2570
box -8 -3 64 105
use XOR2X1  XOR2X1_4
timestamp 1681708930
transform -1 0 1608 0 -1 2570
box -8 -3 64 105
use XOR2X1  XOR2X1_5
timestamp 1681708930
transform -1 0 1664 0 -1 2570
box -8 -3 64 105
use XOR2X1  XOR2X1_6
timestamp 1681708930
transform 1 0 1664 0 -1 2570
box -8 -3 64 105
use FILL  FILL_17
timestamp 1681708930
transform 1 0 1720 0 -1 2570
box -8 -3 16 105
use FILL  FILL_18
timestamp 1681708930
transform 1 0 1728 0 -1 2570
box -8 -3 16 105
use FILL  FILL_19
timestamp 1681708930
transform 1 0 1736 0 -1 2570
box -8 -3 16 105
use FILL  FILL_20
timestamp 1681708930
transform 1 0 1744 0 -1 2570
box -8 -3 16 105
use FILL  FILL_21
timestamp 1681708930
transform 1 0 1752 0 -1 2570
box -8 -3 16 105
use FILL  FILL_22
timestamp 1681708930
transform 1 0 1760 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_0
timestamp 1681708930
transform -1 0 1808 0 -1 2570
box -8 -3 46 105
use INVX2  INVX2_9
timestamp 1681708930
transform 1 0 1808 0 -1 2570
box -9 -3 26 105
use NOR2X1  NOR2X1_0
timestamp 1681708930
transform 1 0 1824 0 -1 2570
box -8 -3 32 105
use FILL  FILL_23
timestamp 1681708930
transform 1 0 1848 0 -1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_0
timestamp 1681708930
transform 1 0 1856 0 -1 2570
box -8 -3 40 105
use INVX2  INVX2_10
timestamp 1681708930
transform 1 0 1888 0 -1 2570
box -9 -3 26 105
use FILL  FILL_24
timestamp 1681708930
transform 1 0 1904 0 -1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_1
timestamp 1681708930
transform 1 0 1912 0 -1 2570
box -8 -3 32 105
use AOI21X1  AOI21X1_0
timestamp 1681708930
transform 1 0 1936 0 -1 2570
box -7 -3 39 105
use FILL  FILL_25
timestamp 1681708930
transform 1 0 1968 0 -1 2570
box -8 -3 16 105
use FILL  FILL_26
timestamp 1681708930
transform 1 0 1976 0 -1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_5
timestamp 1681708930
transform -1 0 2016 0 -1 2570
box -8 -3 34 105
use NAND2X1  NAND2X1_2
timestamp 1681708930
transform 1 0 2016 0 -1 2570
box -8 -3 32 105
use XNOR2X1  XNOR2X1_0
timestamp 1681708930
transform -1 0 2096 0 -1 2570
box -8 -3 64 105
use FILL  FILL_27
timestamp 1681708930
transform 1 0 2096 0 -1 2570
box -8 -3 16 105
use FILL  FILL_28
timestamp 1681708930
transform 1 0 2104 0 -1 2570
box -8 -3 16 105
use XNOR2X1  XNOR2X1_1
timestamp 1681708930
transform -1 0 2168 0 -1 2570
box -8 -3 64 105
use INVX2  INVX2_11
timestamp 1681708930
transform 1 0 2168 0 -1 2570
box -9 -3 26 105
use XNOR2X1  XNOR2X1_2
timestamp 1681708930
transform 1 0 2184 0 -1 2570
box -8 -3 64 105
use FILL  FILL_29
timestamp 1681708930
transform 1 0 2240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_30
timestamp 1681708930
transform 1 0 2248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_31
timestamp 1681708930
transform 1 0 2256 0 -1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_6
timestamp 1681708930
transform 1 0 2264 0 -1 2570
box -8 -3 34 105
use NAND2X1  NAND2X1_3
timestamp 1681708930
transform 1 0 2296 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_4
timestamp 1681708930
transform 1 0 2320 0 -1 2570
box -8 -3 32 105
use NAND3X1  NAND3X1_1
timestamp 1681708930
transform 1 0 2344 0 -1 2570
box -8 -3 40 105
use FILL  FILL_32
timestamp 1681708930
transform 1 0 2376 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_12
timestamp 1681708930
transform 1 0 2384 0 -1 2570
box -9 -3 26 105
use NOR2X1  NOR2X1_2
timestamp 1681708930
transform 1 0 2400 0 -1 2570
box -8 -3 32 105
use AOI22X1  AOI22X1_1
timestamp 1681708930
transform -1 0 2464 0 -1 2570
box -8 -3 46 105
use INVX2  INVX2_13
timestamp 1681708930
transform 1 0 2464 0 -1 2570
box -9 -3 26 105
use NAND3X1  NAND3X1_2
timestamp 1681708930
transform 1 0 2480 0 -1 2570
box -8 -3 40 105
use NOR2X1  NOR2X1_3
timestamp 1681708930
transform -1 0 2536 0 -1 2570
box -8 -3 32 105
use OAI21X1  OAI21X1_7
timestamp 1681708930
transform 1 0 2536 0 -1 2570
box -8 -3 34 105
use FILL  FILL_33
timestamp 1681708930
transform 1 0 2568 0 -1 2570
box -8 -3 16 105
use FILL  FILL_34
timestamp 1681708930
transform 1 0 2576 0 -1 2570
box -8 -3 16 105
use FILL  FILL_35
timestamp 1681708930
transform 1 0 2584 0 -1 2570
box -8 -3 16 105
use FILL  FILL_36
timestamp 1681708930
transform 1 0 2592 0 -1 2570
box -8 -3 16 105
use FILL  FILL_37
timestamp 1681708930
transform 1 0 2600 0 -1 2570
box -8 -3 16 105
use FILL  FILL_38
timestamp 1681708930
transform 1 0 2608 0 -1 2570
box -8 -3 16 105
use FILL  FILL_39
timestamp 1681708930
transform 1 0 2616 0 -1 2570
box -8 -3 16 105
use FILL  FILL_40
timestamp 1681708930
transform 1 0 2624 0 -1 2570
box -8 -3 16 105
use FILL  FILL_41
timestamp 1681708930
transform 1 0 2632 0 -1 2570
box -8 -3 16 105
use FILL  FILL_42
timestamp 1681708930
transform 1 0 2640 0 -1 2570
box -8 -3 16 105
use FILL  FILL_43
timestamp 1681708930
transform 1 0 2648 0 -1 2570
box -8 -3 16 105
use FILL  FILL_44
timestamp 1681708930
transform 1 0 2656 0 -1 2570
box -8 -3 16 105
use top_mod_new_VIA0  top_mod_new_VIA0_3
timestamp 1681708930
transform 1 0 2712 0 1 2470
box -10 -3 10 3
use M3_M2  M3_M2_160
timestamp 1681708930
transform 1 0 100 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_161
timestamp 1681708930
transform 1 0 180 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_162
timestamp 1681708930
transform 1 0 196 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_163
timestamp 1681708930
transform 1 0 212 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_178
timestamp 1681708930
transform 1 0 84 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_179
timestamp 1681708930
transform 1 0 148 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_180
timestamp 1681708930
transform 1 0 188 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_248
timestamp 1681708930
transform 1 0 68 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_207
timestamp 1681708930
transform 1 0 84 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_249
timestamp 1681708930
transform 1 0 100 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_250
timestamp 1681708930
transform 1 0 188 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_225
timestamp 1681708930
transform 1 0 68 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_226
timestamp 1681708930
transform 1 0 148 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_181
timestamp 1681708930
transform 1 0 212 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_182
timestamp 1681708930
transform 1 0 228 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_251
timestamp 1681708930
transform 1 0 220 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_252
timestamp 1681708930
transform 1 0 236 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_227
timestamp 1681708930
transform 1 0 220 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_164
timestamp 1681708930
transform 1 0 268 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_183
timestamp 1681708930
transform 1 0 268 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1681708930
transform 1 0 284 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_253
timestamp 1681708930
transform 1 0 252 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_254
timestamp 1681708930
transform 1 0 276 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_208
timestamp 1681708930
transform 1 0 284 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_165
timestamp 1681708930
transform 1 0 324 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_185
timestamp 1681708930
transform 1 0 308 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_186
timestamp 1681708930
transform 1 0 324 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_255
timestamp 1681708930
transform 1 0 292 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_256
timestamp 1681708930
transform 1 0 300 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_209
timestamp 1681708930
transform 1 0 308 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_257
timestamp 1681708930
transform 1 0 316 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_187
timestamp 1681708930
transform 1 0 356 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_258
timestamp 1681708930
transform 1 0 356 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_166
timestamp 1681708930
transform 1 0 396 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_188
timestamp 1681708930
transform 1 0 380 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_189
timestamp 1681708930
transform 1 0 396 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_210
timestamp 1681708930
transform 1 0 380 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_259
timestamp 1681708930
transform 1 0 388 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_211
timestamp 1681708930
transform 1 0 404 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_167
timestamp 1681708930
transform 1 0 476 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_190
timestamp 1681708930
transform 1 0 452 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_191
timestamp 1681708930
transform 1 0 468 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_192
timestamp 1681708930
transform 1 0 476 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_260
timestamp 1681708930
transform 1 0 436 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_261
timestamp 1681708930
transform 1 0 444 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_212
timestamp 1681708930
transform 1 0 452 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_262
timestamp 1681708930
transform 1 0 476 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_132
timestamp 1681708930
transform 1 0 500 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_168
timestamp 1681708930
transform 1 0 516 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_193
timestamp 1681708930
transform 1 0 484 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_194
timestamp 1681708930
transform 1 0 500 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_195
timestamp 1681708930
transform 1 0 516 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_263
timestamp 1681708930
transform 1 0 492 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_213
timestamp 1681708930
transform 1 0 500 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_264
timestamp 1681708930
transform 1 0 508 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_265
timestamp 1681708930
transform 1 0 548 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_228
timestamp 1681708930
transform 1 0 548 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_196
timestamp 1681708930
transform 1 0 564 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_197
timestamp 1681708930
transform 1 0 580 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_192
timestamp 1681708930
transform 1 0 588 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_266
timestamp 1681708930
transform 1 0 564 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_169
timestamp 1681708930
transform 1 0 628 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_193
timestamp 1681708930
transform 1 0 636 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_198
timestamp 1681708930
transform 1 0 644 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_267
timestamp 1681708930
transform 1 0 612 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_268
timestamp 1681708930
transform 1 0 628 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_269
timestamp 1681708930
transform 1 0 636 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_328
timestamp 1681708930
transform 1 0 620 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_243
timestamp 1681708930
transform 1 0 564 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_244
timestamp 1681708930
transform 1 0 588 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_229
timestamp 1681708930
transform 1 0 628 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_230
timestamp 1681708930
transform 1 0 644 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_245
timestamp 1681708930
transform 1 0 644 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_133
timestamp 1681708930
transform 1 0 716 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_146
timestamp 1681708930
transform 1 0 716 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_151
timestamp 1681708930
transform 1 0 684 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_152
timestamp 1681708930
transform 1 0 700 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_153
timestamp 1681708930
transform 1 0 708 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_199
timestamp 1681708930
transform 1 0 660 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1681708930
transform 1 0 676 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_194
timestamp 1681708930
transform 1 0 684 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_170
timestamp 1681708930
transform 1 0 716 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_154
timestamp 1681708930
transform 1 0 732 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_270
timestamp 1681708930
transform 1 0 676 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_271
timestamp 1681708930
transform 1 0 684 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_214
timestamp 1681708930
transform 1 0 700 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_195
timestamp 1681708930
transform 1 0 732 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_155
timestamp 1681708930
transform 1 0 756 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_201
timestamp 1681708930
transform 1 0 748 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_202
timestamp 1681708930
transform 1 0 764 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_272
timestamp 1681708930
transform 1 0 716 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_273
timestamp 1681708930
transform 1 0 740 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_231
timestamp 1681708930
transform 1 0 668 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_232
timestamp 1681708930
transform 1 0 684 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_246
timestamp 1681708930
transform 1 0 740 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_274
timestamp 1681708930
transform 1 0 764 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_233
timestamp 1681708930
transform 1 0 756 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_247
timestamp 1681708930
transform 1 0 764 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_121
timestamp 1681708930
transform 1 0 828 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_134
timestamp 1681708930
transform 1 0 844 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_156
timestamp 1681708930
transform 1 0 780 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_171
timestamp 1681708930
transform 1 0 788 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_172
timestamp 1681708930
transform 1 0 804 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_173
timestamp 1681708930
transform 1 0 836 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_203
timestamp 1681708930
transform 1 0 788 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_204
timestamp 1681708930
transform 1 0 804 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_205
timestamp 1681708930
transform 1 0 836 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_215
timestamp 1681708930
transform 1 0 780 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_275
timestamp 1681708930
transform 1 0 836 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_276
timestamp 1681708930
transform 1 0 844 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_234
timestamp 1681708930
transform 1 0 836 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_248
timestamp 1681708930
transform 1 0 844 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_122
timestamp 1681708930
transform 1 0 876 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_329
timestamp 1681708930
transform 1 0 868 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_249
timestamp 1681708930
transform 1 0 868 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_157
timestamp 1681708930
transform 1 0 884 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_206
timestamp 1681708930
transform 1 0 884 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_116
timestamp 1681708930
transform 1 0 940 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_123
timestamp 1681708930
transform 1 0 908 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_124
timestamp 1681708930
transform 1 0 940 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_135
timestamp 1681708930
transform 1 0 900 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_207
timestamp 1681708930
transform 1 0 900 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_136
timestamp 1681708930
transform 1 0 972 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_137
timestamp 1681708930
transform 1 0 1020 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_174
timestamp 1681708930
transform 1 0 956 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_175
timestamp 1681708930
transform 1 0 1012 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_196
timestamp 1681708930
transform 1 0 924 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_208
timestamp 1681708930
transform 1 0 972 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_209
timestamp 1681708930
transform 1 0 1004 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_210
timestamp 1681708930
transform 1 0 1012 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_277
timestamp 1681708930
transform 1 0 908 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_278
timestamp 1681708930
transform 1 0 924 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_279
timestamp 1681708930
transform 1 0 1012 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_235
timestamp 1681708930
transform 1 0 972 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_250
timestamp 1681708930
transform 1 0 940 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_251
timestamp 1681708930
transform 1 0 1004 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_158
timestamp 1681708930
transform 1 0 1060 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_280
timestamp 1681708930
transform 1 0 1036 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_281
timestamp 1681708930
transform 1 0 1044 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_236
timestamp 1681708930
transform 1 0 1036 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_252
timestamp 1681708930
transform 1 0 1044 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_176
timestamp 1681708930
transform 1 0 1164 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_197
timestamp 1681708930
transform 1 0 1076 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_138
timestamp 1681708930
transform 1 0 1196 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_211
timestamp 1681708930
transform 1 0 1124 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_212
timestamp 1681708930
transform 1 0 1164 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_213
timestamp 1681708930
transform 1 0 1172 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_282
timestamp 1681708930
transform 1 0 1076 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_216
timestamp 1681708930
transform 1 0 1124 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_283
timestamp 1681708930
transform 1 0 1164 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_217
timestamp 1681708930
transform 1 0 1180 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_159
timestamp 1681708930
transform 1 0 1196 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_177
timestamp 1681708930
transform 1 0 1212 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_198
timestamp 1681708930
transform 1 0 1204 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_284
timestamp 1681708930
transform 1 0 1188 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_285
timestamp 1681708930
transform 1 0 1212 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_286
timestamp 1681708930
transform 1 0 1220 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_125
timestamp 1681708930
transform 1 0 1252 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_139
timestamp 1681708930
transform 1 0 1276 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_178
timestamp 1681708930
transform 1 0 1284 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_160
timestamp 1681708930
transform 1 0 1292 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_214
timestamp 1681708930
transform 1 0 1252 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_215
timestamp 1681708930
transform 1 0 1276 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_199
timestamp 1681708930
transform 1 0 1292 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_287
timestamp 1681708930
transform 1 0 1284 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_161
timestamp 1681708930
transform 1 0 1324 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1681708930
transform 1 0 1316 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_288
timestamp 1681708930
transform 1 0 1308 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_200
timestamp 1681708930
transform 1 0 1324 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_147
timestamp 1681708930
transform 1 0 1372 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_217
timestamp 1681708930
transform 1 0 1372 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_289
timestamp 1681708930
transform 1 0 1340 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_290
timestamp 1681708930
transform 1 0 1348 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_253
timestamp 1681708930
transform 1 0 1340 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_291
timestamp 1681708930
transform 1 0 1396 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_179
timestamp 1681708930
transform 1 0 1420 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_140
timestamp 1681708930
transform 1 0 1452 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_218
timestamp 1681708930
transform 1 0 1428 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_219
timestamp 1681708930
transform 1 0 1452 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_292
timestamp 1681708930
transform 1 0 1420 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_254
timestamp 1681708930
transform 1 0 1412 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_220
timestamp 1681708930
transform 1 0 1492 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_293
timestamp 1681708930
transform 1 0 1476 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_294
timestamp 1681708930
transform 1 0 1484 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_180
timestamp 1681708930
transform 1 0 1572 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_221
timestamp 1681708930
transform 1 0 1548 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_222
timestamp 1681708930
transform 1 0 1572 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_295
timestamp 1681708930
transform 1 0 1540 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1681708930
transform 1 0 1548 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_141
timestamp 1681708930
transform 1 0 1604 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_297
timestamp 1681708930
transform 1 0 1596 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_298
timestamp 1681708930
transform 1 0 1604 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_255
timestamp 1681708930
transform 1 0 1596 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_117
timestamp 1681708930
transform 1 0 1660 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_181
timestamp 1681708930
transform 1 0 1620 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_182
timestamp 1681708930
transform 1 0 1644 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_183
timestamp 1681708930
transform 1 0 1676 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_184
timestamp 1681708930
transform 1 0 1708 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_223
timestamp 1681708930
transform 1 0 1644 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_224
timestamp 1681708930
transform 1 0 1708 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_225
timestamp 1681708930
transform 1 0 1724 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_299
timestamp 1681708930
transform 1 0 1668 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_300
timestamp 1681708930
transform 1 0 1676 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_256
timestamp 1681708930
transform 1 0 1636 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_301
timestamp 1681708930
transform 1 0 1724 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_302
timestamp 1681708930
transform 1 0 1732 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_126
timestamp 1681708930
transform 1 0 1764 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_147
timestamp 1681708930
transform 1 0 1764 0 1 2435
box -2 -2 2 2
use M3_M2  M3_M2_185
timestamp 1681708930
transform 1 0 1756 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_330
timestamp 1681708930
transform 1 0 1756 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_118
timestamp 1681708930
transform 1 0 1780 0 1 2465
box -3 -3 3 3
use M2_M1  M2_M1_162
timestamp 1681708930
transform 1 0 1780 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_186
timestamp 1681708930
transform 1 0 1788 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_127
timestamp 1681708930
transform 1 0 1820 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_142
timestamp 1681708930
transform 1 0 1812 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_148
timestamp 1681708930
transform 1 0 1812 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_163
timestamp 1681708930
transform 1 0 1812 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_187
timestamp 1681708930
transform 1 0 1820 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_226
timestamp 1681708930
transform 1 0 1796 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_227
timestamp 1681708930
transform 1 0 1820 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_303
timestamp 1681708930
transform 1 0 1820 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_119
timestamp 1681708930
transform 1 0 1860 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_143
timestamp 1681708930
transform 1 0 1852 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_149
timestamp 1681708930
transform 1 0 1844 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_164
timestamp 1681708930
transform 1 0 1844 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_228
timestamp 1681708930
transform 1 0 1852 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_304
timestamp 1681708930
transform 1 0 1860 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_165
timestamp 1681708930
transform 1 0 1868 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_229
timestamp 1681708930
transform 1 0 1884 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_305
timestamp 1681708930
transform 1 0 1876 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_218
timestamp 1681708930
transform 1 0 1892 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_331
timestamp 1681708930
transform 1 0 1892 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_306
timestamp 1681708930
transform 1 0 1908 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_120
timestamp 1681708930
transform 1 0 1940 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_128
timestamp 1681708930
transform 1 0 1924 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_150
timestamp 1681708930
transform 1 0 1932 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_144
timestamp 1681708930
transform 1 0 1964 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_145
timestamp 1681708930
transform 1 0 1980 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_148
timestamp 1681708930
transform 1 0 1940 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_166
timestamp 1681708930
transform 1 0 1932 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_188
timestamp 1681708930
transform 1 0 1940 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_167
timestamp 1681708930
transform 1 0 1956 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_168
timestamp 1681708930
transform 1 0 1964 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_230
timestamp 1681708930
transform 1 0 1924 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_307
timestamp 1681708930
transform 1 0 1924 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1681708930
transform 1 0 1940 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1681708930
transform 1 0 1964 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_237
timestamp 1681708930
transform 1 0 1940 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_129
timestamp 1681708930
transform 1 0 2012 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_151
timestamp 1681708930
transform 1 0 2004 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_189
timestamp 1681708930
transform 1 0 1996 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_310
timestamp 1681708930
transform 1 0 1988 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1681708930
transform 1 0 1996 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_238
timestamp 1681708930
transform 1 0 1988 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_152
timestamp 1681708930
transform 1 0 2020 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_169
timestamp 1681708930
transform 1 0 2020 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_146
timestamp 1681708930
transform 1 0 2044 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_153
timestamp 1681708930
transform 1 0 2036 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_170
timestamp 1681708930
transform 1 0 2044 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_231
timestamp 1681708930
transform 1 0 2028 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_257
timestamp 1681708930
transform 1 0 2020 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_232
timestamp 1681708930
transform 1 0 2052 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_233
timestamp 1681708930
transform 1 0 2068 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_312
timestamp 1681708930
transform 1 0 2044 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_313
timestamp 1681708930
transform 1 0 2052 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_258
timestamp 1681708930
transform 1 0 2052 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_154
timestamp 1681708930
transform 1 0 2100 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_171
timestamp 1681708930
transform 1 0 2100 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_234
timestamp 1681708930
transform 1 0 2100 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_219
timestamp 1681708930
transform 1 0 2076 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_314
timestamp 1681708930
transform 1 0 2084 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_220
timestamp 1681708930
transform 1 0 2092 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_235
timestamp 1681708930
transform 1 0 2132 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_221
timestamp 1681708930
transform 1 0 2116 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_315
timestamp 1681708930
transform 1 0 2124 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_332
timestamp 1681708930
transform 1 0 2108 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_259
timestamp 1681708930
transform 1 0 2116 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_155
timestamp 1681708930
transform 1 0 2164 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_201
timestamp 1681708930
transform 1 0 2180 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_236
timestamp 1681708930
transform 1 0 2188 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_316
timestamp 1681708930
transform 1 0 2196 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1681708930
transform 1 0 2244 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_222
timestamp 1681708930
transform 1 0 2252 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_333
timestamp 1681708930
transform 1 0 2252 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_156
timestamp 1681708930
transform 1 0 2284 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_237
timestamp 1681708930
transform 1 0 2268 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_238
timestamp 1681708930
transform 1 0 2300 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1681708930
transform 1 0 2284 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_157
timestamp 1681708930
transform 1 0 2316 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_202
timestamp 1681708930
transform 1 0 2316 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_319
timestamp 1681708930
transform 1 0 2316 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_334
timestamp 1681708930
transform 1 0 2308 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_172
timestamp 1681708930
transform 1 0 2332 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1681708930
transform 1 0 2348 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_239
timestamp 1681708930
transform 1 0 2340 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_173
timestamp 1681708930
transform 1 0 2372 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1681708930
transform 1 0 2372 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_321
timestamp 1681708930
transform 1 0 2380 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_240
timestamp 1681708930
transform 1 0 2380 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_260
timestamp 1681708930
transform 1 0 2372 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_203
timestamp 1681708930
transform 1 0 2436 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_322
timestamp 1681708930
transform 1 0 2428 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_323
timestamp 1681708930
transform 1 0 2436 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_241
timestamp 1681708930
transform 1 0 2452 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_240
timestamp 1681708930
transform 1 0 2476 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_324
timestamp 1681708930
transform 1 0 2468 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_335
timestamp 1681708930
transform 1 0 2460 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_261
timestamp 1681708930
transform 1 0 2460 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_336
timestamp 1681708930
transform 1 0 2476 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_130
timestamp 1681708930
transform 1 0 2492 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_190
timestamp 1681708930
transform 1 0 2500 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_241
timestamp 1681708930
transform 1 0 2492 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_242
timestamp 1681708930
transform 1 0 2500 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_204
timestamp 1681708930
transform 1 0 2516 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_223
timestamp 1681708930
transform 1 0 2500 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_325
timestamp 1681708930
transform 1 0 2508 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_131
timestamp 1681708930
transform 1 0 2532 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_174
timestamp 1681708930
transform 1 0 2532 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_243
timestamp 1681708930
transform 1 0 2532 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_337
timestamp 1681708930
transform 1 0 2524 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_262
timestamp 1681708930
transform 1 0 2524 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_149
timestamp 1681708930
transform 1 0 2548 0 1 2435
box -2 -2 2 2
use M3_M2  M3_M2_191
timestamp 1681708930
transform 1 0 2548 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_175
timestamp 1681708930
transform 1 0 2564 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_176
timestamp 1681708930
transform 1 0 2572 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_244
timestamp 1681708930
transform 1 0 2548 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_263
timestamp 1681708930
transform 1 0 2540 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_205
timestamp 1681708930
transform 1 0 2564 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_150
timestamp 1681708930
transform 1 0 2596 0 1 2435
box -2 -2 2 2
use M3_M2  M3_M2_206
timestamp 1681708930
transform 1 0 2580 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_158
timestamp 1681708930
transform 1 0 2604 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_177
timestamp 1681708930
transform 1 0 2604 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_245
timestamp 1681708930
transform 1 0 2588 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_246
timestamp 1681708930
transform 1 0 2612 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_224
timestamp 1681708930
transform 1 0 2572 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_326
timestamp 1681708930
transform 1 0 2620 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_327
timestamp 1681708930
transform 1 0 2628 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_242
timestamp 1681708930
transform 1 0 2620 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_338
timestamp 1681708930
transform 1 0 2628 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_159
timestamp 1681708930
transform 1 0 2660 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_247
timestamp 1681708930
transform 1 0 2652 0 1 2415
box -2 -2 2 2
use top_mod_new_VIA0  top_mod_new_VIA0_4
timestamp 1681708930
transform 1 0 48 0 1 2370
box -10 -3 10 3
use INVX2  INVX2_14
timestamp 1681708930
transform 1 0 72 0 1 2370
box -9 -3 26 105
use M3_M2  M3_M2_264
timestamp 1681708930
transform 1 0 188 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_8
timestamp 1681708930
transform 1 0 88 0 1 2370
box -8 -3 104 105
use INVX2  INVX2_16
timestamp 1681708930
transform 1 0 184 0 1 2370
box -9 -3 26 105
use OAI22X1  OAI22X1_0
timestamp 1681708930
transform 1 0 200 0 1 2370
box -8 -3 46 105
use INVX2  INVX2_18
timestamp 1681708930
transform -1 0 256 0 1 2370
box -9 -3 26 105
use OAI22X1  OAI22X1_1
timestamp 1681708930
transform 1 0 256 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_2
timestamp 1681708930
transform -1 0 336 0 1 2370
box -8 -3 46 105
use INVX2  INVX2_19
timestamp 1681708930
transform -1 0 352 0 1 2370
box -9 -3 26 105
use FILL  FILL_45
timestamp 1681708930
transform 1 0 352 0 1 2370
box -8 -3 16 105
use FILL  FILL_46
timestamp 1681708930
transform 1 0 360 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_3
timestamp 1681708930
transform -1 0 408 0 1 2370
box -8 -3 46 105
use INVX2  INVX2_20
timestamp 1681708930
transform -1 0 424 0 1 2370
box -9 -3 26 105
use FILL  FILL_47
timestamp 1681708930
transform 1 0 424 0 1 2370
box -8 -3 16 105
use FILL  FILL_48
timestamp 1681708930
transform 1 0 432 0 1 2370
box -8 -3 16 105
use AND2X2  AND2X2_0
timestamp 1681708930
transform 1 0 440 0 1 2370
box -8 -3 40 105
use INVX2  INVX2_21
timestamp 1681708930
transform 1 0 472 0 1 2370
box -9 -3 26 105
use OAI22X1  OAI22X1_4
timestamp 1681708930
transform -1 0 528 0 1 2370
box -8 -3 46 105
use INVX2  INVX2_22
timestamp 1681708930
transform -1 0 544 0 1 2370
box -9 -3 26 105
use FILL  FILL_49
timestamp 1681708930
transform 1 0 544 0 1 2370
box -8 -3 16 105
use FILL  FILL_50
timestamp 1681708930
transform 1 0 552 0 1 2370
box -8 -3 16 105
use XNOR2X1  XNOR2X1_3
timestamp 1681708930
transform -1 0 616 0 1 2370
box -8 -3 64 105
use NOR2X1  NOR2X1_4
timestamp 1681708930
transform 1 0 616 0 1 2370
box -8 -3 32 105
use M3_M2  M3_M2_265
timestamp 1681708930
transform 1 0 652 0 1 2375
box -3 -3 3 3
use FILL  FILL_51
timestamp 1681708930
transform 1 0 640 0 1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_8
timestamp 1681708930
transform 1 0 648 0 1 2370
box -8 -3 34 105
use NAND2X1  NAND2X1_5
timestamp 1681708930
transform 1 0 680 0 1 2370
box -8 -3 32 105
use M3_M2  M3_M2_266
timestamp 1681708930
transform 1 0 716 0 1 2375
box -3 -3 3 3
use NAND3X1  NAND3X1_3
timestamp 1681708930
transform 1 0 704 0 1 2370
box -8 -3 40 105
use NAND2X1  NAND2X1_6
timestamp 1681708930
transform 1 0 736 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_7
timestamp 1681708930
transform 1 0 760 0 1 2370
box -8 -3 32 105
use XNOR2X1  XNOR2X1_4
timestamp 1681708930
transform -1 0 840 0 1 2370
box -8 -3 64 105
use AOI21X1  AOI21X1_1
timestamp 1681708930
transform 1 0 840 0 1 2370
box -7 -3 39 105
use FILL  FILL_61
timestamp 1681708930
transform 1 0 872 0 1 2370
box -8 -3 16 105
use FILL  FILL_62
timestamp 1681708930
transform 1 0 880 0 1 2370
box -8 -3 16 105
use NAND2X1  NAND2X1_8
timestamp 1681708930
transform -1 0 912 0 1 2370
box -8 -3 32 105
use M3_M2  M3_M2_267
timestamp 1681708930
transform 1 0 1012 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_12
timestamp 1681708930
transform 1 0 912 0 1 2370
box -8 -3 104 105
use OAI21X1  OAI21X1_9
timestamp 1681708930
transform 1 0 1008 0 1 2370
box -8 -3 34 105
use NAND2X1  NAND2X1_9
timestamp 1681708930
transform 1 0 1040 0 1 2370
box -8 -3 32 105
use M3_M2  M3_M2_268
timestamp 1681708930
transform 1 0 1164 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_13
timestamp 1681708930
transform 1 0 1064 0 1 2370
box -8 -3 104 105
use OAI21X1  OAI21X1_10
timestamp 1681708930
transform 1 0 1160 0 1 2370
box -8 -3 34 105
use NAND2X1  NAND2X1_10
timestamp 1681708930
transform -1 0 1216 0 1 2370
box -8 -3 32 105
use FILL  FILL_63
timestamp 1681708930
transform 1 0 1216 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_269
timestamp 1681708930
transform 1 0 1284 0 1 2375
box -3 -3 3 3
use XOR2X1  XOR2X1_7
timestamp 1681708930
transform -1 0 1280 0 1 2370
box -8 -3 64 105
use FILL  FILL_64
timestamp 1681708930
transform 1 0 1280 0 1 2370
box -8 -3 16 105
use NAND2X1  NAND2X1_11
timestamp 1681708930
transform -1 0 1312 0 1 2370
box -8 -3 32 105
use FILL  FILL_65
timestamp 1681708930
transform 1 0 1312 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_270
timestamp 1681708930
transform 1 0 1332 0 1 2375
box -3 -3 3 3
use NAND2X1  NAND2X1_12
timestamp 1681708930
transform -1 0 1344 0 1 2370
box -8 -3 32 105
use XOR2X1  XOR2X1_8
timestamp 1681708930
transform -1 0 1400 0 1 2370
box -8 -3 64 105
use FILL  FILL_66
timestamp 1681708930
transform 1 0 1400 0 1 2370
box -8 -3 16 105
use FILL  FILL_67
timestamp 1681708930
transform 1 0 1408 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_271
timestamp 1681708930
transform 1 0 1428 0 1 2375
box -3 -3 3 3
use FILL  FILL_68
timestamp 1681708930
transform 1 0 1416 0 1 2370
box -8 -3 16 105
use XOR2X1  XOR2X1_9
timestamp 1681708930
transform -1 0 1480 0 1 2370
box -8 -3 64 105
use FILL  FILL_69
timestamp 1681708930
transform 1 0 1480 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_272
timestamp 1681708930
transform 1 0 1500 0 1 2375
box -3 -3 3 3
use XNOR2X1  XNOR2X1_5
timestamp 1681708930
transform -1 0 1544 0 1 2370
box -8 -3 64 105
use XOR2X1  XOR2X1_10
timestamp 1681708930
transform -1 0 1600 0 1 2370
box -8 -3 64 105
use FILL  FILL_70
timestamp 1681708930
transform 1 0 1600 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_273
timestamp 1681708930
transform 1 0 1620 0 1 2375
box -3 -3 3 3
use FILL  FILL_71
timestamp 1681708930
transform 1 0 1608 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_274
timestamp 1681708930
transform 1 0 1644 0 1 2375
box -3 -3 3 3
use XOR2X1  XOR2X1_11
timestamp 1681708930
transform -1 0 1672 0 1 2370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_6
timestamp 1681708930
transform 1 0 1672 0 1 2370
box -8 -3 64 105
use FILL  FILL_72
timestamp 1681708930
transform 1 0 1728 0 1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_5
timestamp 1681708930
transform -1 0 1760 0 1 2370
box -8 -3 32 105
use FILL  FILL_73
timestamp 1681708930
transform 1 0 1760 0 1 2370
box -8 -3 16 105
use FILL  FILL_131
timestamp 1681708930
transform 1 0 1768 0 1 2370
box -8 -3 16 105
use FILL  FILL_132
timestamp 1681708930
transform 1 0 1776 0 1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_8
timestamp 1681708930
transform 1 0 1784 0 1 2370
box -8 -3 40 105
use OAI21X1  OAI21X1_13
timestamp 1681708930
transform 1 0 1816 0 1 2370
box -8 -3 34 105
use M3_M2  M3_M2_275
timestamp 1681708930
transform 1 0 1860 0 1 2375
box -3 -3 3 3
use FILL  FILL_133
timestamp 1681708930
transform 1 0 1848 0 1 2370
box -8 -3 16 105
use FILL  FILL_134
timestamp 1681708930
transform 1 0 1856 0 1 2370
box -8 -3 16 105
use FILL  FILL_135
timestamp 1681708930
transform 1 0 1864 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_30
timestamp 1681708930
transform 1 0 1872 0 1 2370
box -9 -3 26 105
use FILL  FILL_137
timestamp 1681708930
transform 1 0 1888 0 1 2370
box -8 -3 16 105
use FILL  FILL_138
timestamp 1681708930
transform 1 0 1896 0 1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_10
timestamp 1681708930
transform 1 0 1904 0 1 2370
box -8 -3 32 105
use NAND3X1  NAND3X1_9
timestamp 1681708930
transform 1 0 1928 0 1 2370
box -8 -3 40 105
use OAI21X1  OAI21X1_14
timestamp 1681708930
transform -1 0 1992 0 1 2370
box -8 -3 34 105
use INVX2  INVX2_31
timestamp 1681708930
transform 1 0 1992 0 1 2370
box -9 -3 26 105
use FILL  FILL_140
timestamp 1681708930
transform 1 0 2008 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_276
timestamp 1681708930
transform 1 0 2028 0 1 2375
box -3 -3 3 3
use FILL  FILL_141
timestamp 1681708930
transform 1 0 2016 0 1 2370
box -8 -3 16 105
use NAND2X1  NAND2X1_15
timestamp 1681708930
transform -1 0 2048 0 1 2370
box -8 -3 32 105
use OAI21X1  OAI21X1_15
timestamp 1681708930
transform -1 0 2080 0 1 2370
box -8 -3 34 105
use NAND2X1  NAND2X1_16
timestamp 1681708930
transform 1 0 2080 0 1 2370
box -8 -3 32 105
use AOI21X1  AOI21X1_4
timestamp 1681708930
transform -1 0 2136 0 1 2370
box -7 -3 39 105
use FILL  FILL_142
timestamp 1681708930
transform 1 0 2136 0 1 2370
box -8 -3 16 105
use FILL  FILL_149
timestamp 1681708930
transform 1 0 2144 0 1 2370
box -8 -3 16 105
use FILL  FILL_151
timestamp 1681708930
transform 1 0 2152 0 1 2370
box -8 -3 16 105
use FILL  FILL_153
timestamp 1681708930
transform 1 0 2160 0 1 2370
box -8 -3 16 105
use FILL  FILL_155
timestamp 1681708930
transform 1 0 2168 0 1 2370
box -8 -3 16 105
use FILL  FILL_157
timestamp 1681708930
transform 1 0 2176 0 1 2370
box -8 -3 16 105
use FILL  FILL_158
timestamp 1681708930
transform 1 0 2184 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_277
timestamp 1681708930
transform 1 0 2244 0 1 2375
box -3 -3 3 3
use XNOR2X1  XNOR2X1_7
timestamp 1681708930
transform -1 0 2248 0 1 2370
box -8 -3 64 105
use NOR2X1  NOR2X1_11
timestamp 1681708930
transform 1 0 2248 0 1 2370
box -8 -3 32 105
use AOI21X1  AOI21X1_6
timestamp 1681708930
transform 1 0 2272 0 1 2370
box -7 -3 39 105
use FILL  FILL_159
timestamp 1681708930
transform 1 0 2304 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_278
timestamp 1681708930
transform 1 0 2348 0 1 2375
box -3 -3 3 3
use NAND2X1  NAND2X1_17
timestamp 1681708930
transform 1 0 2312 0 1 2370
box -8 -3 32 105
use OAI21X1  OAI21X1_17
timestamp 1681708930
transform 1 0 2336 0 1 2370
box -8 -3 34 105
use FILL  FILL_166
timestamp 1681708930
transform 1 0 2368 0 1 2370
box -8 -3 16 105
use XNOR2X1  XNOR2X1_8
timestamp 1681708930
transform 1 0 2376 0 1 2370
box -8 -3 64 105
use AOI21X1  AOI21X1_8
timestamp 1681708930
transform 1 0 2432 0 1 2370
box -7 -3 39 105
use M3_M2  M3_M2_279
timestamp 1681708930
transform 1 0 2484 0 1 2375
box -3 -3 3 3
use FILL  FILL_167
timestamp 1681708930
transform 1 0 2464 0 1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_14
timestamp 1681708930
transform 1 0 2472 0 1 2370
box -8 -3 32 105
use AOI21X1  AOI21X1_9
timestamp 1681708930
transform 1 0 2496 0 1 2370
box -7 -3 39 105
use FILL  FILL_175
timestamp 1681708930
transform 1 0 2528 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_280
timestamp 1681708930
transform 1 0 2564 0 1 2375
box -3 -3 3 3
use NAND3X1  NAND3X1_15
timestamp 1681708930
transform 1 0 2536 0 1 2370
box -8 -3 40 105
use FILL  FILL_176
timestamp 1681708930
transform 1 0 2568 0 1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_16
timestamp 1681708930
transform 1 0 2576 0 1 2370
box -8 -3 40 105
use INVX2  INVX2_35
timestamp 1681708930
transform -1 0 2624 0 1 2370
box -9 -3 26 105
use OR2X1  OR2X1_2
timestamp 1681708930
transform 1 0 2624 0 1 2370
box -8 -3 40 105
use FILL  FILL_177
timestamp 1681708930
transform 1 0 2656 0 1 2370
box -8 -3 16 105
use top_mod_new_VIA0  top_mod_new_VIA0_5
timestamp 1681708930
transform 1 0 2688 0 1 2370
box -10 -3 10 3
use M3_M2  M3_M2_281
timestamp 1681708930
transform 1 0 84 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_309
timestamp 1681708930
transform 1 0 68 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_298
timestamp 1681708930
transform 1 0 164 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_310
timestamp 1681708930
transform 1 0 148 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_353
timestamp 1681708930
transform 1 0 68 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_322
timestamp 1681708930
transform 1 0 84 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_354
timestamp 1681708930
transform 1 0 100 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_413
timestamp 1681708930
transform 1 0 84 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_414
timestamp 1681708930
transform 1 0 148 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_415
timestamp 1681708930
transform 1 0 188 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_299
timestamp 1681708930
transform 1 0 236 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_311
timestamp 1681708930
transform 1 0 220 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_355
timestamp 1681708930
transform 1 0 220 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_356
timestamp 1681708930
transform 1 0 236 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1681708930
transform 1 0 244 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_416
timestamp 1681708930
transform 1 0 212 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_417
timestamp 1681708930
transform 1 0 228 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_358
timestamp 1681708930
transform 1 0 260 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_323
timestamp 1681708930
transform 1 0 276 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_282
timestamp 1681708930
transform 1 0 308 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_324
timestamp 1681708930
transform 1 0 300 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_283
timestamp 1681708930
transform 1 0 356 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_312
timestamp 1681708930
transform 1 0 340 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_300
timestamp 1681708930
transform 1 0 372 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_313
timestamp 1681708930
transform 1 0 396 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_301
timestamp 1681708930
transform 1 0 500 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_314
timestamp 1681708930
transform 1 0 476 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_359
timestamp 1681708930
transform 1 0 324 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_360
timestamp 1681708930
transform 1 0 340 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_361
timestamp 1681708930
transform 1 0 356 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_362
timestamp 1681708930
transform 1 0 372 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_363
timestamp 1681708930
transform 1 0 460 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_418
timestamp 1681708930
transform 1 0 316 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_419
timestamp 1681708930
transform 1 0 332 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_420
timestamp 1681708930
transform 1 0 348 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_344
timestamp 1681708930
transform 1 0 348 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_387
timestamp 1681708930
transform 1 0 340 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_325
timestamp 1681708930
transform 1 0 468 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_364
timestamp 1681708930
transform 1 0 476 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_421
timestamp 1681708930
transform 1 0 396 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_422
timestamp 1681708930
transform 1 0 452 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_423
timestamp 1681708930
transform 1 0 468 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_424
timestamp 1681708930
transform 1 0 484 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_345
timestamp 1681708930
transform 1 0 468 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_388
timestamp 1681708930
transform 1 0 452 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_302
timestamp 1681708930
transform 1 0 524 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_315
timestamp 1681708930
transform 1 0 548 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_365
timestamp 1681708930
transform 1 0 508 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_366
timestamp 1681708930
transform 1 0 524 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_334
timestamp 1681708930
transform 1 0 508 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_425
timestamp 1681708930
transform 1 0 548 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_335
timestamp 1681708930
transform 1 0 572 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_336
timestamp 1681708930
transform 1 0 596 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_284
timestamp 1681708930
transform 1 0 612 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_426
timestamp 1681708930
transform 1 0 604 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_427
timestamp 1681708930
transform 1 0 612 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_358
timestamp 1681708930
transform 1 0 492 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_359
timestamp 1681708930
transform 1 0 516 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_339
timestamp 1681708930
transform 1 0 644 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_367
timestamp 1681708930
transform 1 0 644 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_340
timestamp 1681708930
transform 1 0 700 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_368
timestamp 1681708930
transform 1 0 684 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_369
timestamp 1681708930
transform 1 0 700 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_428
timestamp 1681708930
transform 1 0 668 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_360
timestamp 1681708930
transform 1 0 668 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_370
timestamp 1681708930
transform 1 0 716 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_429
timestamp 1681708930
transform 1 0 700 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_430
timestamp 1681708930
transform 1 0 708 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_346
timestamp 1681708930
transform 1 0 716 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_371
timestamp 1681708930
transform 1 0 740 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_285
timestamp 1681708930
transform 1 0 756 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_286
timestamp 1681708930
transform 1 0 772 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_341
timestamp 1681708930
transform 1 0 756 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_372
timestamp 1681708930
transform 1 0 756 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_373
timestamp 1681708930
transform 1 0 772 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_467
timestamp 1681708930
transform 1 0 764 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_347
timestamp 1681708930
transform 1 0 772 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_287
timestamp 1681708930
transform 1 0 804 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_374
timestamp 1681708930
transform 1 0 796 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_468
timestamp 1681708930
transform 1 0 788 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_361
timestamp 1681708930
transform 1 0 764 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_495
timestamp 1681708930
transform 1 0 772 0 1 2305
box -2 -2 2 2
use M3_M2  M3_M2_377
timestamp 1681708930
transform 1 0 748 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_389
timestamp 1681708930
transform 1 0 764 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_362
timestamp 1681708930
transform 1 0 788 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_378
timestamp 1681708930
transform 1 0 788 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_431
timestamp 1681708930
transform 1 0 812 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_469
timestamp 1681708930
transform 1 0 828 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_288
timestamp 1681708930
transform 1 0 844 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_470
timestamp 1681708930
transform 1 0 836 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_363
timestamp 1681708930
transform 1 0 836 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_375
timestamp 1681708930
transform 1 0 860 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_471
timestamp 1681708930
transform 1 0 868 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_496
timestamp 1681708930
transform 1 0 852 0 1 2305
box -2 -2 2 2
use M3_M2  M3_M2_390
timestamp 1681708930
transform 1 0 844 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_364
timestamp 1681708930
transform 1 0 860 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_376
timestamp 1681708930
transform 1 0 940 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_432
timestamp 1681708930
transform 1 0 908 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_433
timestamp 1681708930
transform 1 0 932 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_472
timestamp 1681708930
transform 1 0 892 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_473
timestamp 1681708930
transform 1 0 900 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_348
timestamp 1681708930
transform 1 0 916 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_474
timestamp 1681708930
transform 1 0 924 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_497
timestamp 1681708930
transform 1 0 884 0 1 2305
box -2 -2 2 2
use M3_M2  M3_M2_379
timestamp 1681708930
transform 1 0 868 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_365
timestamp 1681708930
transform 1 0 900 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_498
timestamp 1681708930
transform 1 0 916 0 1 2305
box -2 -2 2 2
use M3_M2  M3_M2_380
timestamp 1681708930
transform 1 0 908 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_434
timestamp 1681708930
transform 1 0 972 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_326
timestamp 1681708930
transform 1 0 1012 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_327
timestamp 1681708930
transform 1 0 1044 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_435
timestamp 1681708930
transform 1 0 1044 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_475
timestamp 1681708930
transform 1 0 1060 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_377
timestamp 1681708930
transform 1 0 1140 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_366
timestamp 1681708930
transform 1 0 1140 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_378
timestamp 1681708930
transform 1 0 1164 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_303
timestamp 1681708930
transform 1 0 1220 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_436
timestamp 1681708930
transform 1 0 1284 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_316
timestamp 1681708930
transform 1 0 1316 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_379
timestamp 1681708930
transform 1 0 1316 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_476
timestamp 1681708930
transform 1 0 1308 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_289
timestamp 1681708930
transform 1 0 1348 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_317
timestamp 1681708930
transform 1 0 1356 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_380
timestamp 1681708930
transform 1 0 1332 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_328
timestamp 1681708930
transform 1 0 1396 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_381
timestamp 1681708930
transform 1 0 1420 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_437
timestamp 1681708930
transform 1 0 1356 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_438
timestamp 1681708930
transform 1 0 1412 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_337
timestamp 1681708930
transform 1 0 1420 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_342
timestamp 1681708930
transform 1 0 1476 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_382
timestamp 1681708930
transform 1 0 1468 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_439
timestamp 1681708930
transform 1 0 1444 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_349
timestamp 1681708930
transform 1 0 1420 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_350
timestamp 1681708930
transform 1 0 1444 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_391
timestamp 1681708930
transform 1 0 1420 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_367
timestamp 1681708930
transform 1 0 1468 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_318
timestamp 1681708930
transform 1 0 1484 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_343
timestamp 1681708930
transform 1 0 1492 0 1 2345
box -2 -2 2 2
use M3_M2  M3_M2_319
timestamp 1681708930
transform 1 0 1556 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_383
timestamp 1681708930
transform 1 0 1556 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_329
timestamp 1681708930
transform 1 0 1564 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_440
timestamp 1681708930
transform 1 0 1532 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_344
timestamp 1681708930
transform 1 0 1580 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_384
timestamp 1681708930
transform 1 0 1580 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_385
timestamp 1681708930
transform 1 0 1588 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_386
timestamp 1681708930
transform 1 0 1636 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_387
timestamp 1681708930
transform 1 0 1644 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_441
timestamp 1681708930
transform 1 0 1612 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_368
timestamp 1681708930
transform 1 0 1596 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_369
timestamp 1681708930
transform 1 0 1636 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_381
timestamp 1681708930
transform 1 0 1612 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_388
timestamp 1681708930
transform 1 0 1668 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_442
timestamp 1681708930
transform 1 0 1660 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_370
timestamp 1681708930
transform 1 0 1668 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_443
timestamp 1681708930
transform 1 0 1684 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_304
timestamp 1681708930
transform 1 0 1700 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_345
timestamp 1681708930
transform 1 0 1700 0 1 2345
box -2 -2 2 2
use M3_M2  M3_M2_290
timestamp 1681708930
transform 1 0 1740 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_305
timestamp 1681708930
transform 1 0 1732 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_389
timestamp 1681708930
transform 1 0 1724 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_330
timestamp 1681708930
transform 1 0 1732 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_390
timestamp 1681708930
transform 1 0 1740 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_331
timestamp 1681708930
transform 1 0 1748 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_444
timestamp 1681708930
transform 1 0 1724 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_477
timestamp 1681708930
transform 1 0 1732 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_371
timestamp 1681708930
transform 1 0 1732 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_306
timestamp 1681708930
transform 1 0 1764 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_391
timestamp 1681708930
transform 1 0 1772 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_445
timestamp 1681708930
transform 1 0 1764 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_478
timestamp 1681708930
transform 1 0 1756 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_499
timestamp 1681708930
transform 1 0 1748 0 1 2305
box -2 -2 2 2
use M3_M2  M3_M2_291
timestamp 1681708930
transform 1 0 1836 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_320
timestamp 1681708930
transform 1 0 1804 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_321
timestamp 1681708930
transform 1 0 1820 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_346
timestamp 1681708930
transform 1 0 1836 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_392
timestamp 1681708930
transform 1 0 1804 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_393
timestamp 1681708930
transform 1 0 1812 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_394
timestamp 1681708930
transform 1 0 1828 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_446
timestamp 1681708930
transform 1 0 1788 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_447
timestamp 1681708930
transform 1 0 1812 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_448
timestamp 1681708930
transform 1 0 1820 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_372
timestamp 1681708930
transform 1 0 1772 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_382
timestamp 1681708930
transform 1 0 1780 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_479
timestamp 1681708930
transform 1 0 1828 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_347
timestamp 1681708930
transform 1 0 1868 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_449
timestamp 1681708930
transform 1 0 1860 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_338
timestamp 1681708930
transform 1 0 1884 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_348
timestamp 1681708930
transform 1 0 1932 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_395
timestamp 1681708930
transform 1 0 1908 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_396
timestamp 1681708930
transform 1 0 1916 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_450
timestamp 1681708930
transform 1 0 1892 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_451
timestamp 1681708930
transform 1 0 1900 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_332
timestamp 1681708930
transform 1 0 1932 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_339
timestamp 1681708930
transform 1 0 1916 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_452
timestamp 1681708930
transform 1 0 1932 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_453
timestamp 1681708930
transform 1 0 1956 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_349
timestamp 1681708930
transform 1 0 2020 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_454
timestamp 1681708930
transform 1 0 1980 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_455
timestamp 1681708930
transform 1 0 2004 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_480
timestamp 1681708930
transform 1 0 1940 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_481
timestamp 1681708930
transform 1 0 1956 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_482
timestamp 1681708930
transform 1 0 1972 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_392
timestamp 1681708930
transform 1 0 1924 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_351
timestamp 1681708930
transform 1 0 1980 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_483
timestamp 1681708930
transform 1 0 1996 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_500
timestamp 1681708930
transform 1 0 1964 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_501
timestamp 1681708930
transform 1 0 1988 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_397
timestamp 1681708930
transform 1 0 2028 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_333
timestamp 1681708930
transform 1 0 2044 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_398
timestamp 1681708930
transform 1 0 2052 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_456
timestamp 1681708930
transform 1 0 2052 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_457
timestamp 1681708930
transform 1 0 2084 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_352
timestamp 1681708930
transform 1 0 2076 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_484
timestamp 1681708930
transform 1 0 2084 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_393
timestamp 1681708930
transform 1 0 2068 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_458
timestamp 1681708930
transform 1 0 2100 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_502
timestamp 1681708930
transform 1 0 2108 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_485
timestamp 1681708930
transform 1 0 2124 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_292
timestamp 1681708930
transform 1 0 2172 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_293
timestamp 1681708930
transform 1 0 2196 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_307
timestamp 1681708930
transform 1 0 2204 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_350
timestamp 1681708930
transform 1 0 2204 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_399
timestamp 1681708930
transform 1 0 2188 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_400
timestamp 1681708930
transform 1 0 2204 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_459
timestamp 1681708930
transform 1 0 2180 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_353
timestamp 1681708930
transform 1 0 2180 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_294
timestamp 1681708930
transform 1 0 2244 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_308
timestamp 1681708930
transform 1 0 2236 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_351
timestamp 1681708930
transform 1 0 2244 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_401
timestamp 1681708930
transform 1 0 2236 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_402
timestamp 1681708930
transform 1 0 2244 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_403
timestamp 1681708930
transform 1 0 2260 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_460
timestamp 1681708930
transform 1 0 2212 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_461
timestamp 1681708930
transform 1 0 2220 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_373
timestamp 1681708930
transform 1 0 2212 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_383
timestamp 1681708930
transform 1 0 2188 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_340
timestamp 1681708930
transform 1 0 2260 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_486
timestamp 1681708930
transform 1 0 2236 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_354
timestamp 1681708930
transform 1 0 2244 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_404
timestamp 1681708930
transform 1 0 2284 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_462
timestamp 1681708930
transform 1 0 2276 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_355
timestamp 1681708930
transform 1 0 2276 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_356
timestamp 1681708930
transform 1 0 2300 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_295
timestamp 1681708930
transform 1 0 2340 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_405
timestamp 1681708930
transform 1 0 2332 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_463
timestamp 1681708930
transform 1 0 2324 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_352
timestamp 1681708930
transform 1 0 2348 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_406
timestamp 1681708930
transform 1 0 2356 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_407
timestamp 1681708930
transform 1 0 2372 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_341
timestamp 1681708930
transform 1 0 2364 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_487
timestamp 1681708930
transform 1 0 2364 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_503
timestamp 1681708930
transform 1 0 2364 0 1 2305
box -2 -2 2 2
use M3_M2  M3_M2_384
timestamp 1681708930
transform 1 0 2364 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_488
timestamp 1681708930
transform 1 0 2412 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_296
timestamp 1681708930
transform 1 0 2436 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_504
timestamp 1681708930
transform 1 0 2420 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_505
timestamp 1681708930
transform 1 0 2428 0 1 2305
box -2 -2 2 2
use M3_M2  M3_M2_374
timestamp 1681708930
transform 1 0 2436 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_385
timestamp 1681708930
transform 1 0 2420 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_464
timestamp 1681708930
transform 1 0 2452 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_386
timestamp 1681708930
transform 1 0 2452 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_297
timestamp 1681708930
transform 1 0 2476 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_408
timestamp 1681708930
transform 1 0 2468 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_342
timestamp 1681708930
transform 1 0 2468 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_489
timestamp 1681708930
transform 1 0 2468 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_409
timestamp 1681708930
transform 1 0 2500 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_410
timestamp 1681708930
transform 1 0 2540 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_465
timestamp 1681708930
transform 1 0 2524 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_490
timestamp 1681708930
transform 1 0 2500 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_491
timestamp 1681708930
transform 1 0 2508 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_357
timestamp 1681708930
transform 1 0 2516 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_492
timestamp 1681708930
transform 1 0 2532 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_493
timestamp 1681708930
transform 1 0 2556 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_506
timestamp 1681708930
transform 1 0 2516 0 1 2305
box -2 -2 2 2
use M3_M2  M3_M2_375
timestamp 1681708930
transform 1 0 2524 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_376
timestamp 1681708930
transform 1 0 2556 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_411
timestamp 1681708930
transform 1 0 2588 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_343
timestamp 1681708930
transform 1 0 2588 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_494
timestamp 1681708930
transform 1 0 2580 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_507
timestamp 1681708930
transform 1 0 2564 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_412
timestamp 1681708930
transform 1 0 2652 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_466
timestamp 1681708930
transform 1 0 2668 0 1 2325
box -2 -2 2 2
use top_mod_new_VIA0  top_mod_new_VIA0_6
timestamp 1681708930
transform 1 0 24 0 1 2270
box -10 -3 10 3
use INVX2  INVX2_15
timestamp 1681708930
transform 1 0 72 0 -1 2370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_9
timestamp 1681708930
transform 1 0 88 0 -1 2370
box -8 -3 104 105
use INVX2  INVX2_17
timestamp 1681708930
transform 1 0 184 0 -1 2370
box -9 -3 26 105
use OAI22X1  OAI22X1_5
timestamp 1681708930
transform 1 0 200 0 -1 2370
box -8 -3 46 105
use M3_M2  M3_M2_394
timestamp 1681708930
transform 1 0 252 0 1 2275
box -3 -3 3 3
use FILL  FILL_52
timestamp 1681708930
transform 1 0 240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_53
timestamp 1681708930
transform 1 0 248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_54
timestamp 1681708930
transform 1 0 256 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_23
timestamp 1681708930
transform 1 0 264 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_24
timestamp 1681708930
transform 1 0 280 0 -1 2370
box -9 -3 26 105
use FILL  FILL_55
timestamp 1681708930
transform 1 0 296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_56
timestamp 1681708930
transform 1 0 304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_57
timestamp 1681708930
transform 1 0 312 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_6
timestamp 1681708930
transform 1 0 320 0 -1 2370
box -8 -3 46 105
use M3_M2  M3_M2_395
timestamp 1681708930
transform 1 0 428 0 1 2275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_10
timestamp 1681708930
transform 1 0 360 0 -1 2370
box -8 -3 104 105
use OAI22X1  OAI22X1_7
timestamp 1681708930
transform -1 0 496 0 -1 2370
box -8 -3 46 105
use INVX2  INVX2_25
timestamp 1681708930
transform -1 0 512 0 -1 2370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_11
timestamp 1681708930
transform 1 0 512 0 -1 2370
box -8 -3 104 105
use FILL  FILL_58
timestamp 1681708930
transform 1 0 608 0 -1 2370
box -8 -3 16 105
use FILL  FILL_59
timestamp 1681708930
transform 1 0 616 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_26
timestamp 1681708930
transform -1 0 640 0 -1 2370
box -9 -3 26 105
use FILL  FILL_60
timestamp 1681708930
transform 1 0 640 0 -1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_6
timestamp 1681708930
transform 1 0 648 0 -1 2370
box -8 -3 32 105
use AOI21X1  AOI21X1_2
timestamp 1681708930
transform 1 0 672 0 -1 2370
box -7 -3 39 105
use FILL  FILL_74
timestamp 1681708930
transform 1 0 704 0 -1 2370
box -8 -3 16 105
use FILL  FILL_75
timestamp 1681708930
transform 1 0 712 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_27
timestamp 1681708930
transform 1 0 720 0 -1 2370
box -9 -3 26 105
use NOR2X1  NOR2X1_7
timestamp 1681708930
transform -1 0 760 0 -1 2370
box -8 -3 32 105
use M3_M2  M3_M2_396
timestamp 1681708930
transform 1 0 780 0 1 2275
box -3 -3 3 3
use NAND3X1  NAND3X1_4
timestamp 1681708930
transform 1 0 760 0 -1 2370
box -8 -3 40 105
use M3_M2  M3_M2_397
timestamp 1681708930
transform 1 0 804 0 1 2275
box -3 -3 3 3
use FILL  FILL_76
timestamp 1681708930
transform 1 0 792 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_11
timestamp 1681708930
transform 1 0 800 0 -1 2370
box -8 -3 34 105
use FILL  FILL_77
timestamp 1681708930
transform 1 0 832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_78
timestamp 1681708930
transform 1 0 840 0 -1 2370
box -8 -3 16 105
use FILL  FILL_79
timestamp 1681708930
transform 1 0 848 0 -1 2370
box -8 -3 16 105
use FILL  FILL_80
timestamp 1681708930
transform 1 0 856 0 -1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_5
timestamp 1681708930
transform 1 0 864 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_6
timestamp 1681708930
transform 1 0 896 0 -1 2370
box -8 -3 40 105
use INVX2  INVX2_28
timestamp 1681708930
transform -1 0 944 0 -1 2370
box -9 -3 26 105
use FILL  FILL_81
timestamp 1681708930
transform 1 0 944 0 -1 2370
box -8 -3 16 105
use FILL  FILL_82
timestamp 1681708930
transform 1 0 952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_83
timestamp 1681708930
transform 1 0 960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_84
timestamp 1681708930
transform 1 0 968 0 -1 2370
box -8 -3 16 105
use FILL  FILL_85
timestamp 1681708930
transform 1 0 976 0 -1 2370
box -8 -3 16 105
use FILL  FILL_86
timestamp 1681708930
transform 1 0 984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_87
timestamp 1681708930
transform 1 0 992 0 -1 2370
box -8 -3 16 105
use FILL  FILL_88
timestamp 1681708930
transform 1 0 1000 0 -1 2370
box -8 -3 16 105
use FILL  FILL_89
timestamp 1681708930
transform 1 0 1008 0 -1 2370
box -8 -3 16 105
use FILL  FILL_90
timestamp 1681708930
transform 1 0 1016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_91
timestamp 1681708930
transform 1 0 1024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_92
timestamp 1681708930
transform 1 0 1032 0 -1 2370
box -8 -3 16 105
use FILL  FILL_93
timestamp 1681708930
transform 1 0 1040 0 -1 2370
box -8 -3 16 105
use FILL  FILL_94
timestamp 1681708930
transform 1 0 1048 0 -1 2370
box -8 -3 16 105
use FILL  FILL_95
timestamp 1681708930
transform 1 0 1056 0 -1 2370
box -8 -3 16 105
use FILL  FILL_96
timestamp 1681708930
transform 1 0 1064 0 -1 2370
box -8 -3 16 105
use NAND2X1  NAND2X1_13
timestamp 1681708930
transform -1 0 1096 0 -1 2370
box -8 -3 32 105
use FILL  FILL_97
timestamp 1681708930
transform 1 0 1096 0 -1 2370
box -8 -3 16 105
use FILL  FILL_98
timestamp 1681708930
transform 1 0 1104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_99
timestamp 1681708930
transform 1 0 1112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_100
timestamp 1681708930
transform 1 0 1120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_101
timestamp 1681708930
transform 1 0 1128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_102
timestamp 1681708930
transform 1 0 1136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_103
timestamp 1681708930
transform 1 0 1144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_104
timestamp 1681708930
transform 1 0 1152 0 -1 2370
box -8 -3 16 105
use FILL  FILL_105
timestamp 1681708930
transform 1 0 1160 0 -1 2370
box -8 -3 16 105
use FILL  FILL_106
timestamp 1681708930
transform 1 0 1168 0 -1 2370
box -8 -3 16 105
use FILL  FILL_107
timestamp 1681708930
transform 1 0 1176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_108
timestamp 1681708930
transform 1 0 1184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_109
timestamp 1681708930
transform 1 0 1192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_110
timestamp 1681708930
transform 1 0 1200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_111
timestamp 1681708930
transform 1 0 1208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_112
timestamp 1681708930
transform 1 0 1216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_113
timestamp 1681708930
transform 1 0 1224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_114
timestamp 1681708930
transform 1 0 1232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_115
timestamp 1681708930
transform 1 0 1240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_116
timestamp 1681708930
transform 1 0 1248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_117
timestamp 1681708930
transform 1 0 1256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_118
timestamp 1681708930
transform 1 0 1264 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_12
timestamp 1681708930
transform 1 0 1272 0 -1 2370
box -8 -3 34 105
use FILL  FILL_119
timestamp 1681708930
transform 1 0 1304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_120
timestamp 1681708930
transform 1 0 1312 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_14
timestamp 1681708930
transform 1 0 1320 0 -1 2370
box -8 -3 104 105
use XOR2X1  XOR2X1_12
timestamp 1681708930
transform -1 0 1472 0 -1 2370
box -8 -3 64 105
use FILL  FILL_121
timestamp 1681708930
transform 1 0 1472 0 -1 2370
box -8 -3 16 105
use FILL  FILL_122
timestamp 1681708930
transform 1 0 1480 0 -1 2370
box -8 -3 16 105
use FILL  FILL_123
timestamp 1681708930
transform 1 0 1488 0 -1 2370
box -8 -3 16 105
use FILL  FILL_124
timestamp 1681708930
transform 1 0 1496 0 -1 2370
box -8 -3 16 105
use XOR2X1  XOR2X1_13
timestamp 1681708930
transform 1 0 1504 0 -1 2370
box -8 -3 64 105
use M3_M2  M3_M2_398
timestamp 1681708930
transform 1 0 1588 0 1 2275
box -3 -3 3 3
use NOR2X1  NOR2X1_8
timestamp 1681708930
transform -1 0 1584 0 -1 2370
box -8 -3 32 105
use XOR2X1  XOR2X1_14
timestamp 1681708930
transform -1 0 1640 0 -1 2370
box -8 -3 64 105
use FILL  FILL_125
timestamp 1681708930
transform 1 0 1640 0 -1 2370
box -8 -3 16 105
use FILL  FILL_126
timestamp 1681708930
transform 1 0 1648 0 -1 2370
box -8 -3 16 105
use FILL  FILL_127
timestamp 1681708930
transform 1 0 1656 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_29
timestamp 1681708930
transform 1 0 1664 0 -1 2370
box -9 -3 26 105
use FILL  FILL_128
timestamp 1681708930
transform 1 0 1680 0 -1 2370
box -8 -3 16 105
use FILL  FILL_129
timestamp 1681708930
transform 1 0 1688 0 -1 2370
box -8 -3 16 105
use AOI21X1  AOI21X1_3
timestamp 1681708930
transform -1 0 1728 0 -1 2370
box -7 -3 39 105
use NAND3X1  NAND3X1_7
timestamp 1681708930
transform 1 0 1728 0 -1 2370
box -8 -3 40 105
use FILL  FILL_130
timestamp 1681708930
transform 1 0 1760 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_2
timestamp 1681708930
transform 1 0 1768 0 -1 2370
box -8 -3 46 105
use NAND2X1  NAND2X1_14
timestamp 1681708930
transform 1 0 1808 0 -1 2370
box -8 -3 32 105
use OR2X1  OR2X1_0
timestamp 1681708930
transform 1 0 1832 0 -1 2370
box -8 -3 40 105
use FILL  FILL_136
timestamp 1681708930
transform 1 0 1864 0 -1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_9
timestamp 1681708930
transform 1 0 1872 0 -1 2370
box -8 -3 32 105
use FILL  FILL_139
timestamp 1681708930
transform 1 0 1896 0 -1 2370
box -8 -3 16 105
use AOI21X1  AOI21X1_5
timestamp 1681708930
transform 1 0 1904 0 -1 2370
box -7 -3 39 105
use NAND3X1  NAND3X1_10
timestamp 1681708930
transform -1 0 1968 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_11
timestamp 1681708930
transform 1 0 1968 0 -1 2370
box -8 -3 40 105
use INVX2  INVX2_32
timestamp 1681708930
transform -1 0 2016 0 -1 2370
box -9 -3 26 105
use OR2X1  OR2X1_1
timestamp 1681708930
transform 1 0 2016 0 -1 2370
box -8 -3 40 105
use FILL  FILL_143
timestamp 1681708930
transform 1 0 2048 0 -1 2370
box -8 -3 16 105
use FILL  FILL_144
timestamp 1681708930
transform 1 0 2056 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_33
timestamp 1681708930
transform 1 0 2064 0 -1 2370
box -9 -3 26 105
use FILL  FILL_145
timestamp 1681708930
transform 1 0 2080 0 -1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_12
timestamp 1681708930
transform 1 0 2088 0 -1 2370
box -8 -3 40 105
use FILL  FILL_146
timestamp 1681708930
transform 1 0 2120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_147
timestamp 1681708930
transform 1 0 2128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_148
timestamp 1681708930
transform 1 0 2136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_150
timestamp 1681708930
transform 1 0 2144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_152
timestamp 1681708930
transform 1 0 2152 0 -1 2370
box -8 -3 16 105
use FILL  FILL_154
timestamp 1681708930
transform 1 0 2160 0 -1 2370
box -8 -3 16 105
use FILL  FILL_156
timestamp 1681708930
transform 1 0 2168 0 -1 2370
box -8 -3 16 105
use AOI21X1  AOI21X1_7
timestamp 1681708930
transform 1 0 2176 0 -1 2370
box -7 -3 39 105
use OAI21X1  OAI21X1_16
timestamp 1681708930
transform 1 0 2208 0 -1 2370
box -8 -3 34 105
use NOR2X1  NOR2X1_12
timestamp 1681708930
transform 1 0 2240 0 -1 2370
box -8 -3 32 105
use FILL  FILL_160
timestamp 1681708930
transform 1 0 2264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_161
timestamp 1681708930
transform 1 0 2272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_162
timestamp 1681708930
transform 1 0 2280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_163
timestamp 1681708930
transform 1 0 2288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_164
timestamp 1681708930
transform 1 0 2296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_165
timestamp 1681708930
transform 1 0 2304 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_34
timestamp 1681708930
transform 1 0 2312 0 -1 2370
box -9 -3 26 105
use NOR2X1  NOR2X1_13
timestamp 1681708930
transform -1 0 2352 0 -1 2370
box -8 -3 32 105
use FILL  FILL_168
timestamp 1681708930
transform 1 0 2352 0 -1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_13
timestamp 1681708930
transform 1 0 2360 0 -1 2370
box -8 -3 40 105
use FILL  FILL_169
timestamp 1681708930
transform 1 0 2392 0 -1 2370
box -8 -3 16 105
use FILL  FILL_170
timestamp 1681708930
transform 1 0 2400 0 -1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_14
timestamp 1681708930
transform 1 0 2408 0 -1 2370
box -8 -3 40 105
use FILL  FILL_171
timestamp 1681708930
transform 1 0 2440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_172
timestamp 1681708930
transform 1 0 2448 0 -1 2370
box -8 -3 16 105
use FILL  FILL_173
timestamp 1681708930
transform 1 0 2456 0 -1 2370
box -8 -3 16 105
use FILL  FILL_174
timestamp 1681708930
transform 1 0 2464 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_18
timestamp 1681708930
transform 1 0 2472 0 -1 2370
box -8 -3 34 105
use NAND3X1  NAND3X1_17
timestamp 1681708930
transform -1 0 2536 0 -1 2370
box -8 -3 40 105
use INVX2  INVX2_36
timestamp 1681708930
transform 1 0 2536 0 -1 2370
box -9 -3 26 105
use NAND3X1  NAND3X1_18
timestamp 1681708930
transform 1 0 2552 0 -1 2370
box -8 -3 40 105
use FILL  FILL_178
timestamp 1681708930
transform 1 0 2584 0 -1 2370
box -8 -3 16 105
use XOR2X1  XOR2X1_15
timestamp 1681708930
transform 1 0 2592 0 -1 2370
box -8 -3 64 105
use FILL  FILL_179
timestamp 1681708930
transform 1 0 2648 0 -1 2370
box -8 -3 16 105
use FILL  FILL_180
timestamp 1681708930
transform 1 0 2656 0 -1 2370
box -8 -3 16 105
use top_mod_new_VIA0  top_mod_new_VIA0_7
timestamp 1681708930
transform 1 0 2712 0 1 2270
box -10 -3 10 3
use M2_M1  M2_M1_536
timestamp 1681708930
transform 1 0 76 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_603
timestamp 1681708930
transform 1 0 68 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_604
timestamp 1681708930
transform 1 0 92 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_500
timestamp 1681708930
transform 1 0 68 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_430
timestamp 1681708930
transform 1 0 108 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_399
timestamp 1681708930
transform 1 0 188 0 1 2265
box -3 -3 3 3
use M2_M1  M2_M1_537
timestamp 1681708930
transform 1 0 108 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_538
timestamp 1681708930
transform 1 0 116 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_539
timestamp 1681708930
transform 1 0 172 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_431
timestamp 1681708930
transform 1 0 220 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_432
timestamp 1681708930
transform 1 0 236 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_540
timestamp 1681708930
transform 1 0 220 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_541
timestamp 1681708930
transform 1 0 236 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_451
timestamp 1681708930
transform 1 0 244 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_605
timestamp 1681708930
transform 1 0 196 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_606
timestamp 1681708930
transform 1 0 212 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_607
timestamp 1681708930
transform 1 0 228 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_608
timestamp 1681708930
transform 1 0 244 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_475
timestamp 1681708930
transform 1 0 172 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_476
timestamp 1681708930
transform 1 0 228 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_407
timestamp 1681708930
transform 1 0 260 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_609
timestamp 1681708930
transform 1 0 260 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_477
timestamp 1681708930
transform 1 0 260 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_501
timestamp 1681708930
transform 1 0 260 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_417
timestamp 1681708930
transform 1 0 284 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_542
timestamp 1681708930
transform 1 0 284 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_610
timestamp 1681708930
transform 1 0 284 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_408
timestamp 1681708930
transform 1 0 300 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_433
timestamp 1681708930
transform 1 0 316 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_543
timestamp 1681708930
transform 1 0 316 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_544
timestamp 1681708930
transform 1 0 324 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_409
timestamp 1681708930
transform 1 0 348 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_545
timestamp 1681708930
transform 1 0 340 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_611
timestamp 1681708930
transform 1 0 348 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_478
timestamp 1681708930
transform 1 0 348 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_502
timestamp 1681708930
transform 1 0 340 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_434
timestamp 1681708930
transform 1 0 364 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_435
timestamp 1681708930
transform 1 0 380 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_546
timestamp 1681708930
transform 1 0 364 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_452
timestamp 1681708930
transform 1 0 372 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_547
timestamp 1681708930
transform 1 0 380 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_612
timestamp 1681708930
transform 1 0 372 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_613
timestamp 1681708930
transform 1 0 412 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_614
timestamp 1681708930
transform 1 0 420 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_503
timestamp 1681708930
transform 1 0 420 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_418
timestamp 1681708930
transform 1 0 460 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_548
timestamp 1681708930
transform 1 0 444 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_615
timestamp 1681708930
transform 1 0 452 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_479
timestamp 1681708930
transform 1 0 444 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_549
timestamp 1681708930
transform 1 0 468 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_550
timestamp 1681708930
transform 1 0 484 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_480
timestamp 1681708930
transform 1 0 468 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_616
timestamp 1681708930
transform 1 0 492 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_504
timestamp 1681708930
transform 1 0 492 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_436
timestamp 1681708930
transform 1 0 532 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_551
timestamp 1681708930
transform 1 0 516 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_552
timestamp 1681708930
transform 1 0 532 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_617
timestamp 1681708930
transform 1 0 524 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_553
timestamp 1681708930
transform 1 0 588 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_618
timestamp 1681708930
transform 1 0 580 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_619
timestamp 1681708930
transform 1 0 588 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_481
timestamp 1681708930
transform 1 0 580 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_482
timestamp 1681708930
transform 1 0 604 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_410
timestamp 1681708930
transform 1 0 628 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_419
timestamp 1681708930
transform 1 0 628 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_437
timestamp 1681708930
transform 1 0 636 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_554
timestamp 1681708930
transform 1 0 612 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_555
timestamp 1681708930
transform 1 0 620 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_556
timestamp 1681708930
transform 1 0 636 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_557
timestamp 1681708930
transform 1 0 660 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_620
timestamp 1681708930
transform 1 0 644 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_621
timestamp 1681708930
transform 1 0 660 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_420
timestamp 1681708930
transform 1 0 668 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_438
timestamp 1681708930
transform 1 0 676 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_558
timestamp 1681708930
transform 1 0 668 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_559
timestamp 1681708930
transform 1 0 676 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_622
timestamp 1681708930
transform 1 0 684 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_403
timestamp 1681708930
transform 1 0 700 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_411
timestamp 1681708930
transform 1 0 700 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_514
timestamp 1681708930
transform 1 0 724 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_671
timestamp 1681708930
transform 1 0 732 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_623
timestamp 1681708930
transform 1 0 772 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_483
timestamp 1681708930
transform 1 0 772 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_400
timestamp 1681708930
transform 1 0 812 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_421
timestamp 1681708930
transform 1 0 804 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_422
timestamp 1681708930
transform 1 0 828 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_560
timestamp 1681708930
transform 1 0 788 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_561
timestamp 1681708930
transform 1 0 796 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_453
timestamp 1681708930
transform 1 0 812 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_562
timestamp 1681708930
transform 1 0 828 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_624
timestamp 1681708930
transform 1 0 796 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_625
timestamp 1681708930
transform 1 0 804 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_505
timestamp 1681708930
transform 1 0 788 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_672
timestamp 1681708930
transform 1 0 820 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_404
timestamp 1681708930
transform 1 0 844 0 1 2255
box -3 -3 3 3
use M2_M1  M2_M1_508
timestamp 1681708930
transform 1 0 844 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_515
timestamp 1681708930
transform 1 0 844 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_454
timestamp 1681708930
transform 1 0 844 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_563
timestamp 1681708930
transform 1 0 852 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_564
timestamp 1681708930
transform 1 0 868 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_405
timestamp 1681708930
transform 1 0 892 0 1 2255
box -3 -3 3 3
use M2_M1  M2_M1_626
timestamp 1681708930
transform 1 0 908 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_423
timestamp 1681708930
transform 1 0 932 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_516
timestamp 1681708930
transform 1 0 932 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_517
timestamp 1681708930
transform 1 0 940 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_455
timestamp 1681708930
transform 1 0 932 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_565
timestamp 1681708930
transform 1 0 956 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_464
timestamp 1681708930
transform 1 0 956 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_627
timestamp 1681708930
transform 1 0 964 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_628
timestamp 1681708930
transform 1 0 980 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_673
timestamp 1681708930
transform 1 0 972 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_484
timestamp 1681708930
transform 1 0 980 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_566
timestamp 1681708930
transform 1 0 1012 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_567
timestamp 1681708930
transform 1 0 1020 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_629
timestamp 1681708930
transform 1 0 1004 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_465
timestamp 1681708930
transform 1 0 1020 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_485
timestamp 1681708930
transform 1 0 1012 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_518
timestamp 1681708930
transform 1 0 1044 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_439
timestamp 1681708930
transform 1 0 1060 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_568
timestamp 1681708930
transform 1 0 1084 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_569
timestamp 1681708930
transform 1 0 1140 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_456
timestamp 1681708930
transform 1 0 1148 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_519
timestamp 1681708930
transform 1 0 1172 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_570
timestamp 1681708930
transform 1 0 1156 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_630
timestamp 1681708930
transform 1 0 1044 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_631
timestamp 1681708930
transform 1 0 1060 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_466
timestamp 1681708930
transform 1 0 1140 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_632
timestamp 1681708930
transform 1 0 1148 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_486
timestamp 1681708930
transform 1 0 1044 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_487
timestamp 1681708930
transform 1 0 1084 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_440
timestamp 1681708930
transform 1 0 1228 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_441
timestamp 1681708930
transform 1 0 1260 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_571
timestamp 1681708930
transform 1 0 1180 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_572
timestamp 1681708930
transform 1 0 1212 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_457
timestamp 1681708930
transform 1 0 1236 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_633
timestamp 1681708930
transform 1 0 1172 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_467
timestamp 1681708930
transform 1 0 1212 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_520
timestamp 1681708930
transform 1 0 1308 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_573
timestamp 1681708930
transform 1 0 1284 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_634
timestamp 1681708930
transform 1 0 1260 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_635
timestamp 1681708930
transform 1 0 1276 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_488
timestamp 1681708930
transform 1 0 1172 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_489
timestamp 1681708930
transform 1 0 1212 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_458
timestamp 1681708930
transform 1 0 1308 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_636
timestamp 1681708930
transform 1 0 1308 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_468
timestamp 1681708930
transform 1 0 1316 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_442
timestamp 1681708930
transform 1 0 1340 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_574
timestamp 1681708930
transform 1 0 1364 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_575
timestamp 1681708930
transform 1 0 1420 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_637
timestamp 1681708930
transform 1 0 1324 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_638
timestamp 1681708930
transform 1 0 1340 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_469
timestamp 1681708930
transform 1 0 1364 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_521
timestamp 1681708930
transform 1 0 1460 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_401
timestamp 1681708930
transform 1 0 1476 0 1 2265
box -3 -3 3 3
use M2_M1  M2_M1_509
timestamp 1681708930
transform 1 0 1484 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_510
timestamp 1681708930
transform 1 0 1500 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_522
timestamp 1681708930
transform 1 0 1492 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_576
timestamp 1681708930
transform 1 0 1484 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_639
timestamp 1681708930
transform 1 0 1500 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_490
timestamp 1681708930
transform 1 0 1500 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_577
timestamp 1681708930
transform 1 0 1524 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_424
timestamp 1681708930
transform 1 0 1540 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_402
timestamp 1681708930
transform 1 0 1564 0 1 2265
box -3 -3 3 3
use M2_M1  M2_M1_578
timestamp 1681708930
transform 1 0 1548 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_579
timestamp 1681708930
transform 1 0 1564 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_425
timestamp 1681708930
transform 1 0 1588 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_580
timestamp 1681708930
transform 1 0 1588 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_640
timestamp 1681708930
transform 1 0 1564 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_641
timestamp 1681708930
transform 1 0 1572 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_642
timestamp 1681708930
transform 1 0 1596 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_491
timestamp 1681708930
transform 1 0 1572 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_674
timestamp 1681708930
transform 1 0 1588 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_581
timestamp 1681708930
transform 1 0 1652 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_643
timestamp 1681708930
transform 1 0 1644 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_492
timestamp 1681708930
transform 1 0 1644 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_644
timestamp 1681708930
transform 1 0 1660 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_470
timestamp 1681708930
transform 1 0 1668 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_523
timestamp 1681708930
transform 1 0 1692 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_645
timestamp 1681708930
transform 1 0 1700 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_524
timestamp 1681708930
transform 1 0 1716 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_582
timestamp 1681708930
transform 1 0 1716 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_583
timestamp 1681708930
transform 1 0 1724 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_471
timestamp 1681708930
transform 1 0 1716 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_646
timestamp 1681708930
transform 1 0 1748 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_675
timestamp 1681708930
transform 1 0 1740 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_493
timestamp 1681708930
transform 1 0 1748 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_584
timestamp 1681708930
transform 1 0 1764 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_494
timestamp 1681708930
transform 1 0 1764 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_585
timestamp 1681708930
transform 1 0 1772 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_647
timestamp 1681708930
transform 1 0 1772 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_459
timestamp 1681708930
transform 1 0 1788 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_586
timestamp 1681708930
transform 1 0 1796 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_460
timestamp 1681708930
transform 1 0 1804 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_587
timestamp 1681708930
transform 1 0 1812 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_648
timestamp 1681708930
transform 1 0 1788 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_649
timestamp 1681708930
transform 1 0 1804 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_472
timestamp 1681708930
transform 1 0 1820 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_650
timestamp 1681708930
transform 1 0 1828 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_495
timestamp 1681708930
transform 1 0 1804 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_496
timestamp 1681708930
transform 1 0 1836 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_525
timestamp 1681708930
transform 1 0 1844 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_511
timestamp 1681708930
transform 1 0 1860 0 1 2235
box -2 -2 2 2
use M3_M2  M3_M2_443
timestamp 1681708930
transform 1 0 1876 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_406
timestamp 1681708930
transform 1 0 1948 0 1 2255
box -3 -3 3 3
use M2_M1  M2_M1_526
timestamp 1681708930
transform 1 0 1884 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_473
timestamp 1681708930
transform 1 0 1860 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_444
timestamp 1681708930
transform 1 0 1908 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_445
timestamp 1681708930
transform 1 0 1924 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_588
timestamp 1681708930
transform 1 0 1908 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_651
timestamp 1681708930
transform 1 0 1868 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_652
timestamp 1681708930
transform 1 0 1892 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_497
timestamp 1681708930
transform 1 0 1868 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_446
timestamp 1681708930
transform 1 0 1972 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_589
timestamp 1681708930
transform 1 0 1972 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_653
timestamp 1681708930
transform 1 0 1940 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_654
timestamp 1681708930
transform 1 0 1948 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_506
timestamp 1681708930
transform 1 0 1892 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_507
timestamp 1681708930
transform 1 0 1908 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_508
timestamp 1681708930
transform 1 0 1924 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_655
timestamp 1681708930
transform 1 0 1996 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_656
timestamp 1681708930
transform 1 0 2004 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_509
timestamp 1681708930
transform 1 0 1980 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_590
timestamp 1681708930
transform 1 0 2060 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_657
timestamp 1681708930
transform 1 0 2052 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_658
timestamp 1681708930
transform 1 0 2068 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_447
timestamp 1681708930
transform 1 0 2100 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_591
timestamp 1681708930
transform 1 0 2100 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_659
timestamp 1681708930
transform 1 0 2124 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_510
timestamp 1681708930
transform 1 0 2100 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_660
timestamp 1681708930
transform 1 0 2188 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_511
timestamp 1681708930
transform 1 0 2188 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_412
timestamp 1681708930
transform 1 0 2212 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_527
timestamp 1681708930
transform 1 0 2212 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_592
timestamp 1681708930
transform 1 0 2212 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_593
timestamp 1681708930
transform 1 0 2220 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_594
timestamp 1681708930
transform 1 0 2228 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_413
timestamp 1681708930
transform 1 0 2252 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_528
timestamp 1681708930
transform 1 0 2252 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_661
timestamp 1681708930
transform 1 0 2228 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_662
timestamp 1681708930
transform 1 0 2236 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_474
timestamp 1681708930
transform 1 0 2244 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_498
timestamp 1681708930
transform 1 0 2228 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_461
timestamp 1681708930
transform 1 0 2276 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_663
timestamp 1681708930
transform 1 0 2316 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_664
timestamp 1681708930
transform 1 0 2324 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_512
timestamp 1681708930
transform 1 0 2292 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_499
timestamp 1681708930
transform 1 0 2324 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_414
timestamp 1681708930
transform 1 0 2364 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_426
timestamp 1681708930
transform 1 0 2356 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_448
timestamp 1681708930
transform 1 0 2356 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_427
timestamp 1681708930
transform 1 0 2388 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_529
timestamp 1681708930
transform 1 0 2380 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_595
timestamp 1681708930
transform 1 0 2356 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_596
timestamp 1681708930
transform 1 0 2364 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_665
timestamp 1681708930
transform 1 0 2348 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_676
timestamp 1681708930
transform 1 0 2340 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_462
timestamp 1681708930
transform 1 0 2372 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_597
timestamp 1681708930
transform 1 0 2380 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_535
timestamp 1681708930
transform 1 0 2388 0 1 2217
box -2 -2 2 2
use M2_M1  M2_M1_598
timestamp 1681708930
transform 1 0 2412 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_666
timestamp 1681708930
transform 1 0 2388 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_677
timestamp 1681708930
transform 1 0 2412 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_415
timestamp 1681708930
transform 1 0 2452 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_416
timestamp 1681708930
transform 1 0 2508 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_512
timestamp 1681708930
transform 1 0 2460 0 1 2235
box -2 -2 2 2
use M3_M2  M3_M2_428
timestamp 1681708930
transform 1 0 2476 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_513
timestamp 1681708930
transform 1 0 2500 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_530
timestamp 1681708930
transform 1 0 2452 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_449
timestamp 1681708930
transform 1 0 2460 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_531
timestamp 1681708930
transform 1 0 2476 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_532
timestamp 1681708930
transform 1 0 2500 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_533
timestamp 1681708930
transform 1 0 2508 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_534
timestamp 1681708930
transform 1 0 2524 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_599
timestamp 1681708930
transform 1 0 2492 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_463
timestamp 1681708930
transform 1 0 2500 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_667
timestamp 1681708930
transform 1 0 2484 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_450
timestamp 1681708930
transform 1 0 2564 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_429
timestamp 1681708930
transform 1 0 2588 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_600
timestamp 1681708930
transform 1 0 2564 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_601
timestamp 1681708930
transform 1 0 2580 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1681708930
transform 1 0 2532 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_513
timestamp 1681708930
transform 1 0 2564 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_602
timestamp 1681708930
transform 1 0 2596 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_669
timestamp 1681708930
transform 1 0 2588 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_670
timestamp 1681708930
transform 1 0 2660 0 1 2205
box -2 -2 2 2
use top_mod_new_VIA0  top_mod_new_VIA0_8
timestamp 1681708930
transform 1 0 48 0 1 2170
box -10 -3 10 3
use INVX2  INVX2_37
timestamp 1681708930
transform 1 0 72 0 1 2170
box -9 -3 26 105
use M3_M2  M3_M2_514
timestamp 1681708930
transform 1 0 116 0 1 2175
box -3 -3 3 3
use INVX2  INVX2_39
timestamp 1681708930
transform 1 0 88 0 1 2170
box -9 -3 26 105
use FILL  FILL_181
timestamp 1681708930
transform 1 0 104 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_515
timestamp 1681708930
transform 1 0 164 0 1 2175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_15
timestamp 1681708930
transform -1 0 208 0 1 2170
box -8 -3 104 105
use M3_M2  M3_M2_516
timestamp 1681708930
transform 1 0 252 0 1 2175
box -3 -3 3 3
use OAI22X1  OAI22X1_8
timestamp 1681708930
transform -1 0 248 0 1 2170
box -8 -3 46 105
use FILL  FILL_182
timestamp 1681708930
transform 1 0 248 0 1 2170
box -8 -3 16 105
use FILL  FILL_183
timestamp 1681708930
transform 1 0 256 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_40
timestamp 1681708930
transform 1 0 264 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_41
timestamp 1681708930
transform 1 0 280 0 1 2170
box -9 -3 26 105
use FILL  FILL_184
timestamp 1681708930
transform 1 0 296 0 1 2170
box -8 -3 16 105
use FILL  FILL_200
timestamp 1681708930
transform 1 0 304 0 1 2170
box -8 -3 16 105
use FILL  FILL_202
timestamp 1681708930
transform 1 0 312 0 1 2170
box -8 -3 16 105
use FILL  FILL_204
timestamp 1681708930
transform 1 0 320 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_43
timestamp 1681708930
transform -1 0 344 0 1 2170
box -9 -3 26 105
use FILL  FILL_205
timestamp 1681708930
transform 1 0 344 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_517
timestamp 1681708930
transform 1 0 396 0 1 2175
box -3 -3 3 3
use OAI22X1  OAI22X1_11
timestamp 1681708930
transform -1 0 392 0 1 2170
box -8 -3 46 105
use FILL  FILL_206
timestamp 1681708930
transform 1 0 392 0 1 2170
box -8 -3 16 105
use FILL  FILL_207
timestamp 1681708930
transform 1 0 400 0 1 2170
box -8 -3 16 105
use FILL  FILL_208
timestamp 1681708930
transform 1 0 408 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_44
timestamp 1681708930
transform 1 0 416 0 1 2170
box -9 -3 26 105
use M3_M2  M3_M2_518
timestamp 1681708930
transform 1 0 452 0 1 2175
box -3 -3 3 3
use INVX2  INVX2_45
timestamp 1681708930
transform 1 0 432 0 1 2170
box -9 -3 26 105
use FILL  FILL_209
timestamp 1681708930
transform 1 0 448 0 1 2170
box -8 -3 16 105
use AND2X2  AND2X2_1
timestamp 1681708930
transform 1 0 456 0 1 2170
box -8 -3 40 105
use FILL  FILL_215
timestamp 1681708930
transform 1 0 488 0 1 2170
box -8 -3 16 105
use FILL  FILL_216
timestamp 1681708930
transform 1 0 496 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_12
timestamp 1681708930
transform -1 0 544 0 1 2170
box -8 -3 46 105
use FILL  FILL_217
timestamp 1681708930
transform 1 0 544 0 1 2170
box -8 -3 16 105
use FILL  FILL_218
timestamp 1681708930
transform 1 0 552 0 1 2170
box -8 -3 16 105
use FILL  FILL_219
timestamp 1681708930
transform 1 0 560 0 1 2170
box -8 -3 16 105
use FILL  FILL_220
timestamp 1681708930
transform 1 0 568 0 1 2170
box -8 -3 16 105
use FILL  FILL_221
timestamp 1681708930
transform 1 0 576 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_46
timestamp 1681708930
transform 1 0 584 0 1 2170
box -9 -3 26 105
use FILL  FILL_222
timestamp 1681708930
transform 1 0 600 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_519
timestamp 1681708930
transform 1 0 620 0 1 2175
box -3 -3 3 3
use FILL  FILL_223
timestamp 1681708930
transform 1 0 608 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_3
timestamp 1681708930
transform 1 0 616 0 1 2170
box -8 -3 46 105
use INVX2  INVX2_47
timestamp 1681708930
transform 1 0 656 0 1 2170
box -9 -3 26 105
use FILL  FILL_224
timestamp 1681708930
transform 1 0 672 0 1 2170
box -8 -3 16 105
use FILL  FILL_225
timestamp 1681708930
transform 1 0 680 0 1 2170
box -8 -3 16 105
use FILL  FILL_226
timestamp 1681708930
transform 1 0 688 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_520
timestamp 1681708930
transform 1 0 716 0 1 2175
box -3 -3 3 3
use OAI21X1  OAI21X1_19
timestamp 1681708930
transform 1 0 696 0 1 2170
box -8 -3 34 105
use FILL  FILL_227
timestamp 1681708930
transform 1 0 728 0 1 2170
box -8 -3 16 105
use FILL  FILL_228
timestamp 1681708930
transform 1 0 736 0 1 2170
box -8 -3 16 105
use FILL  FILL_229
timestamp 1681708930
transform 1 0 744 0 1 2170
box -8 -3 16 105
use FILL  FILL_230
timestamp 1681708930
transform 1 0 752 0 1 2170
box -8 -3 16 105
use FILL  FILL_231
timestamp 1681708930
transform 1 0 760 0 1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_15
timestamp 1681708930
transform 1 0 768 0 1 2170
box -8 -3 32 105
use AOI21X1  AOI21X1_10
timestamp 1681708930
transform 1 0 792 0 1 2170
box -7 -3 39 105
use INVX2  INVX2_48
timestamp 1681708930
transform 1 0 824 0 1 2170
box -9 -3 26 105
use FILL  FILL_232
timestamp 1681708930
transform 1 0 840 0 1 2170
box -8 -3 16 105
use FILL  FILL_244
timestamp 1681708930
transform 1 0 848 0 1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_20
timestamp 1681708930
transform 1 0 856 0 1 2170
box -8 -3 40 105
use FILL  FILL_245
timestamp 1681708930
transform 1 0 888 0 1 2170
box -8 -3 16 105
use FILL  FILL_246
timestamp 1681708930
transform 1 0 896 0 1 2170
box -8 -3 16 105
use FILL  FILL_247
timestamp 1681708930
transform 1 0 904 0 1 2170
box -8 -3 16 105
use FILL  FILL_248
timestamp 1681708930
transform 1 0 912 0 1 2170
box -8 -3 16 105
use FILL  FILL_249
timestamp 1681708930
transform 1 0 920 0 1 2170
box -8 -3 16 105
use FILL  FILL_250
timestamp 1681708930
transform 1 0 928 0 1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_21
timestamp 1681708930
transform -1 0 968 0 1 2170
box -8 -3 34 105
use OR2X1  OR2X1_3
timestamp 1681708930
transform 1 0 968 0 1 2170
box -8 -3 40 105
use FILL  FILL_251
timestamp 1681708930
transform 1 0 1000 0 1 2170
box -8 -3 16 105
use FILL  FILL_252
timestamp 1681708930
transform 1 0 1008 0 1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_22
timestamp 1681708930
transform 1 0 1016 0 1 2170
box -8 -3 34 105
use M3_M2  M3_M2_521
timestamp 1681708930
transform 1 0 1148 0 1 2175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_18
timestamp 1681708930
transform 1 0 1048 0 1 2170
box -8 -3 104 105
use OAI21X1  OAI21X1_23
timestamp 1681708930
transform 1 0 1144 0 1 2170
box -8 -3 34 105
use M3_M2  M3_M2_522
timestamp 1681708930
transform 1 0 1276 0 1 2175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_19
timestamp 1681708930
transform -1 0 1272 0 1 2170
box -8 -3 104 105
use OAI21X1  OAI21X1_24
timestamp 1681708930
transform 1 0 1272 0 1 2170
box -8 -3 34 105
use NAND2X1  NAND2X1_18
timestamp 1681708930
transform -1 0 1328 0 1 2170
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_20
timestamp 1681708930
transform 1 0 1328 0 1 2170
box -8 -3 104 105
use FILL  FILL_253
timestamp 1681708930
transform 1 0 1424 0 1 2170
box -8 -3 16 105
use FILL  FILL_254
timestamp 1681708930
transform 1 0 1432 0 1 2170
box -8 -3 16 105
use FILL  FILL_255
timestamp 1681708930
transform 1 0 1440 0 1 2170
box -8 -3 16 105
use FILL  FILL_256
timestamp 1681708930
transform 1 0 1448 0 1 2170
box -8 -3 16 105
use FILL  FILL_257
timestamp 1681708930
transform 1 0 1456 0 1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_21
timestamp 1681708930
transform -1 0 1496 0 1 2170
box -8 -3 40 105
use FILL  FILL_258
timestamp 1681708930
transform 1 0 1496 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_523
timestamp 1681708930
transform 1 0 1532 0 1 2175
box -3 -3 3 3
use INVX2  INVX2_51
timestamp 1681708930
transform 1 0 1504 0 1 2170
box -9 -3 26 105
use FILL  FILL_259
timestamp 1681708930
transform 1 0 1520 0 1 2170
box -8 -3 16 105
use FILL  FILL_260
timestamp 1681708930
transform 1 0 1528 0 1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_19
timestamp 1681708930
transform -1 0 1560 0 1 2170
box -8 -3 32 105
use AOI21X1  AOI21X1_11
timestamp 1681708930
transform 1 0 1560 0 1 2170
box -7 -3 39 105
use XOR2X1  XOR2X1_18
timestamp 1681708930
transform 1 0 1592 0 1 2170
box -8 -3 64 105
use FILL  FILL_261
timestamp 1681708930
transform 1 0 1648 0 1 2170
box -8 -3 16 105
use FILL  FILL_262
timestamp 1681708930
transform 1 0 1656 0 1 2170
box -8 -3 16 105
use FILL  FILL_263
timestamp 1681708930
transform 1 0 1664 0 1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_20
timestamp 1681708930
transform 1 0 1672 0 1 2170
box -8 -3 32 105
use FILL  FILL_264
timestamp 1681708930
transform 1 0 1696 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_524
timestamp 1681708930
transform 1 0 1716 0 1 2175
box -3 -3 3 3
use FILL  FILL_265
timestamp 1681708930
transform 1 0 1704 0 1 2170
box -8 -3 16 105
use FILL  FILL_266
timestamp 1681708930
transform 1 0 1712 0 1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_16
timestamp 1681708930
transform -1 0 1744 0 1 2170
box -8 -3 32 105
use M3_M2  M3_M2_525
timestamp 1681708930
transform 1 0 1764 0 1 2175
box -3 -3 3 3
use INVX2  INVX2_52
timestamp 1681708930
transform 1 0 1744 0 1 2170
box -9 -3 26 105
use FILL  FILL_267
timestamp 1681708930
transform 1 0 1760 0 1 2170
box -8 -3 16 105
use FILL  FILL_268
timestamp 1681708930
transform 1 0 1768 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_4
timestamp 1681708930
transform 1 0 1776 0 1 2170
box -8 -3 46 105
use INVX2  INVX2_53
timestamp 1681708930
transform -1 0 1832 0 1 2170
box -9 -3 26 105
use FILL  FILL_269
timestamp 1681708930
transform 1 0 1832 0 1 2170
box -8 -3 16 105
use FILL  FILL_270
timestamp 1681708930
transform 1 0 1840 0 1 2170
box -8 -3 16 105
use FILL  FILL_271
timestamp 1681708930
transform 1 0 1848 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_526
timestamp 1681708930
transform 1 0 1876 0 1 2175
box -3 -3 3 3
use NAND3X1  NAND3X1_24
timestamp 1681708930
transform 1 0 1856 0 1 2170
box -8 -3 40 105
use XOR2X1  XOR2X1_23
timestamp 1681708930
transform -1 0 1944 0 1 2170
box -8 -3 64 105
use M3_M2  M3_M2_527
timestamp 1681708930
transform 1 0 2004 0 1 2175
box -3 -3 3 3
use XOR2X1  XOR2X1_24
timestamp 1681708930
transform -1 0 2000 0 1 2170
box -8 -3 64 105
use M3_M2  M3_M2_528
timestamp 1681708930
transform 1 0 2044 0 1 2175
box -3 -3 3 3
use XOR2X1  XOR2X1_25
timestamp 1681708930
transform 1 0 2000 0 1 2170
box -8 -3 64 105
use FILL  FILL_287
timestamp 1681708930
transform 1 0 2056 0 1 2170
box -8 -3 16 105
use FILL  FILL_288
timestamp 1681708930
transform 1 0 2064 0 1 2170
box -8 -3 16 105
use XOR2X1  XOR2X1_26
timestamp 1681708930
transform 1 0 2072 0 1 2170
box -8 -3 64 105
use FILL  FILL_289
timestamp 1681708930
transform 1 0 2128 0 1 2170
box -8 -3 16 105
use FILL  FILL_290
timestamp 1681708930
transform 1 0 2136 0 1 2170
box -8 -3 16 105
use FILL  FILL_291
timestamp 1681708930
transform 1 0 2144 0 1 2170
box -8 -3 16 105
use FILL  FILL_292
timestamp 1681708930
transform 1 0 2152 0 1 2170
box -8 -3 16 105
use FILL  FILL_293
timestamp 1681708930
transform 1 0 2160 0 1 2170
box -8 -3 16 105
use FILL  FILL_294
timestamp 1681708930
transform 1 0 2168 0 1 2170
box -8 -3 16 105
use FILL  FILL_295
timestamp 1681708930
transform 1 0 2176 0 1 2170
box -8 -3 16 105
use FILL  FILL_302
timestamp 1681708930
transform 1 0 2184 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_57
timestamp 1681708930
transform 1 0 2192 0 1 2170
box -9 -3 26 105
use NAND2X1  NAND2X1_24
timestamp 1681708930
transform -1 0 2232 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_25
timestamp 1681708930
transform 1 0 2232 0 1 2170
box -8 -3 32 105
use XNOR2X1  XNOR2X1_9
timestamp 1681708930
transform 1 0 2256 0 1 2170
box -8 -3 64 105
use AOI21X1  AOI21X1_12
timestamp 1681708930
transform 1 0 2312 0 1 2170
box -7 -3 39 105
use FILL  FILL_304
timestamp 1681708930
transform 1 0 2344 0 1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_29
timestamp 1681708930
transform 1 0 2352 0 1 2170
box -8 -3 34 105
use AOI21X1  AOI21X1_13
timestamp 1681708930
transform 1 0 2384 0 1 2170
box -7 -3 39 105
use FILL  FILL_308
timestamp 1681708930
transform 1 0 2416 0 1 2170
box -8 -3 16 105
use FILL  FILL_309
timestamp 1681708930
transform 1 0 2424 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_59
timestamp 1681708930
transform 1 0 2432 0 1 2170
box -9 -3 26 105
use NAND3X1  NAND3X1_28
timestamp 1681708930
transform 1 0 2448 0 1 2170
box -8 -3 40 105
use INVX2  INVX2_60
timestamp 1681708930
transform 1 0 2480 0 1 2170
box -9 -3 26 105
use NAND3X1  NAND3X1_29
timestamp 1681708930
transform 1 0 2496 0 1 2170
box -8 -3 40 105
use XOR2X1  XOR2X1_31
timestamp 1681708930
transform 1 0 2528 0 1 2170
box -8 -3 64 105
use FILL  FILL_310
timestamp 1681708930
transform 1 0 2584 0 1 2170
box -8 -3 16 105
use FILL  FILL_311
timestamp 1681708930
transform 1 0 2592 0 1 2170
box -8 -3 16 105
use XOR2X1  XOR2X1_32
timestamp 1681708930
transform -1 0 2656 0 1 2170
box -8 -3 64 105
use FILL  FILL_312
timestamp 1681708930
transform 1 0 2656 0 1 2170
box -8 -3 16 105
use top_mod_new_VIA0  top_mod_new_VIA0_9
timestamp 1681708930
transform 1 0 2688 0 1 2170
box -10 -3 10 3
use M2_M1  M2_M1_684
timestamp 1681708930
transform 1 0 68 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_618
timestamp 1681708930
transform 1 0 68 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_582
timestamp 1681708930
transform 1 0 92 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_598
timestamp 1681708930
transform 1 0 140 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_569
timestamp 1681708930
transform 1 0 180 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_570
timestamp 1681708930
transform 1 0 212 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_685
timestamp 1681708930
transform 1 0 180 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_686
timestamp 1681708930
transform 1 0 196 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_756
timestamp 1681708930
transform 1 0 172 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_757
timestamp 1681708930
transform 1 0 188 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_599
timestamp 1681708930
transform 1 0 196 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_758
timestamp 1681708930
transform 1 0 212 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_619
timestamp 1681708930
transform 1 0 212 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_687
timestamp 1681708930
transform 1 0 236 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_600
timestamp 1681708930
transform 1 0 236 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_759
timestamp 1681708930
transform 1 0 244 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_620
timestamp 1681708930
transform 1 0 228 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_643
timestamp 1681708930
transform 1 0 236 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_541
timestamp 1681708930
transform 1 0 284 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_688
timestamp 1681708930
transform 1 0 252 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_689
timestamp 1681708930
transform 1 0 260 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_690
timestamp 1681708930
transform 1 0 276 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_760
timestamp 1681708930
transform 1 0 252 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_601
timestamp 1681708930
transform 1 0 260 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_761
timestamp 1681708930
transform 1 0 268 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_762
timestamp 1681708930
transform 1 0 284 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_621
timestamp 1681708930
transform 1 0 284 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_644
timestamp 1681708930
transform 1 0 292 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_665
timestamp 1681708930
transform 1 0 308 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_763
timestamp 1681708930
transform 1 0 324 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_571
timestamp 1681708930
transform 1 0 348 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_529
timestamp 1681708930
transform 1 0 436 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_691
timestamp 1681708930
transform 1 0 364 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_583
timestamp 1681708930
transform 1 0 412 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_530
timestamp 1681708930
transform 1 0 452 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_679
timestamp 1681708930
transform 1 0 452 0 1 2145
box -2 -2 2 2
use M3_M2  M3_M2_584
timestamp 1681708930
transform 1 0 452 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_764
timestamp 1681708930
transform 1 0 388 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_765
timestamp 1681708930
transform 1 0 444 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_766
timestamp 1681708930
transform 1 0 452 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_622
timestamp 1681708930
transform 1 0 388 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_645
timestamp 1681708930
transform 1 0 356 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_666
timestamp 1681708930
transform 1 0 372 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_542
timestamp 1681708930
transform 1 0 460 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_692
timestamp 1681708930
transform 1 0 484 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_767
timestamp 1681708930
transform 1 0 484 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_623
timestamp 1681708930
transform 1 0 484 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_667
timestamp 1681708930
transform 1 0 492 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_585
timestamp 1681708930
transform 1 0 524 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_531
timestamp 1681708930
transform 1 0 628 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_543
timestamp 1681708930
transform 1 0 612 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_693
timestamp 1681708930
transform 1 0 540 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_586
timestamp 1681708930
transform 1 0 564 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_532
timestamp 1681708930
transform 1 0 676 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_544
timestamp 1681708930
transform 1 0 644 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_545
timestamp 1681708930
transform 1 0 660 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_694
timestamp 1681708930
transform 1 0 628 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_768
timestamp 1681708930
transform 1 0 564 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_602
timestamp 1681708930
transform 1 0 588 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_546
timestamp 1681708930
transform 1 0 692 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_695
timestamp 1681708930
transform 1 0 676 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_587
timestamp 1681708930
transform 1 0 700 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_696
timestamp 1681708930
transform 1 0 716 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_769
timestamp 1681708930
transform 1 0 620 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_603
timestamp 1681708930
transform 1 0 644 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_770
timestamp 1681708930
transform 1 0 652 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_604
timestamp 1681708930
transform 1 0 684 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_771
timestamp 1681708930
transform 1 0 692 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_605
timestamp 1681708930
transform 1 0 700 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_772
timestamp 1681708930
transform 1 0 716 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_624
timestamp 1681708930
transform 1 0 628 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_606
timestamp 1681708930
transform 1 0 740 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_625
timestamp 1681708930
transform 1 0 676 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_815
timestamp 1681708930
transform 1 0 684 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_626
timestamp 1681708930
transform 1 0 692 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_816
timestamp 1681708930
transform 1 0 708 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_627
timestamp 1681708930
transform 1 0 716 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_834
timestamp 1681708930
transform 1 0 684 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_654
timestamp 1681708930
transform 1 0 652 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_655
timestamp 1681708930
transform 1 0 684 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_697
timestamp 1681708930
transform 1 0 772 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_698
timestamp 1681708930
transform 1 0 788 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_773
timestamp 1681708930
transform 1 0 780 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_607
timestamp 1681708930
transform 1 0 788 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_817
timestamp 1681708930
transform 1 0 812 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_668
timestamp 1681708930
transform 1 0 796 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_699
timestamp 1681708930
transform 1 0 836 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_533
timestamp 1681708930
transform 1 0 940 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_700
timestamp 1681708930
transform 1 0 860 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_534
timestamp 1681708930
transform 1 0 956 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_701
timestamp 1681708930
transform 1 0 956 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_774
timestamp 1681708930
transform 1 0 908 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_775
timestamp 1681708930
transform 1 0 940 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_776
timestamp 1681708930
transform 1 0 948 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_818
timestamp 1681708930
transform 1 0 972 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_547
timestamp 1681708930
transform 1 0 996 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_548
timestamp 1681708930
transform 1 0 1060 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_702
timestamp 1681708930
transform 1 0 996 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_588
timestamp 1681708930
transform 1 0 1044 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_589
timestamp 1681708930
transform 1 0 1076 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_703
timestamp 1681708930
transform 1 0 1084 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_777
timestamp 1681708930
transform 1 0 1044 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_778
timestamp 1681708930
transform 1 0 1076 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_628
timestamp 1681708930
transform 1 0 1044 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_704
timestamp 1681708930
transform 1 0 1108 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_705
timestamp 1681708930
transform 1 0 1116 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_779
timestamp 1681708930
transform 1 0 1100 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_819
timestamp 1681708930
transform 1 0 1084 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_608
timestamp 1681708930
transform 1 0 1108 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_706
timestamp 1681708930
transform 1 0 1164 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_780
timestamp 1681708930
transform 1 0 1140 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_669
timestamp 1681708930
transform 1 0 1140 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_707
timestamp 1681708930
transform 1 0 1204 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_781
timestamp 1681708930
transform 1 0 1188 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_782
timestamp 1681708930
transform 1 0 1196 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_820
timestamp 1681708930
transform 1 0 1188 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_656
timestamp 1681708930
transform 1 0 1188 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_609
timestamp 1681708930
transform 1 0 1204 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_670
timestamp 1681708930
transform 1 0 1212 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_708
timestamp 1681708930
transform 1 0 1244 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_821
timestamp 1681708930
transform 1 0 1244 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_657
timestamp 1681708930
transform 1 0 1244 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_549
timestamp 1681708930
transform 1 0 1284 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_709
timestamp 1681708930
transform 1 0 1276 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_710
timestamp 1681708930
transform 1 0 1284 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_646
timestamp 1681708930
transform 1 0 1268 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_658
timestamp 1681708930
transform 1 0 1276 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_550
timestamp 1681708930
transform 1 0 1332 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_711
timestamp 1681708930
transform 1 0 1332 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_712
timestamp 1681708930
transform 1 0 1340 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_783
timestamp 1681708930
transform 1 0 1300 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_659
timestamp 1681708930
transform 1 0 1308 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_551
timestamp 1681708930
transform 1 0 1388 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_552
timestamp 1681708930
transform 1 0 1420 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_713
timestamp 1681708930
transform 1 0 1388 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_714
timestamp 1681708930
transform 1 0 1396 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_784
timestamp 1681708930
transform 1 0 1364 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_535
timestamp 1681708930
transform 1 0 1500 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_572
timestamp 1681708930
transform 1 0 1484 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_715
timestamp 1681708930
transform 1 0 1444 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_716
timestamp 1681708930
transform 1 0 1460 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_785
timestamp 1681708930
transform 1 0 1420 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_786
timestamp 1681708930
transform 1 0 1452 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_647
timestamp 1681708930
transform 1 0 1396 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_671
timestamp 1681708930
transform 1 0 1420 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_553
timestamp 1681708930
transform 1 0 1508 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_554
timestamp 1681708930
transform 1 0 1564 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_680
timestamp 1681708930
transform 1 0 1564 0 1 2145
box -2 -2 2 2
use M3_M2  M3_M2_573
timestamp 1681708930
transform 1 0 1572 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_717
timestamp 1681708930
transform 1 0 1508 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_718
timestamp 1681708930
transform 1 0 1524 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_590
timestamp 1681708930
transform 1 0 1540 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_719
timestamp 1681708930
transform 1 0 1556 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_787
timestamp 1681708930
transform 1 0 1500 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_788
timestamp 1681708930
transform 1 0 1516 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_789
timestamp 1681708930
transform 1 0 1532 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_790
timestamp 1681708930
transform 1 0 1540 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_822
timestamp 1681708930
transform 1 0 1468 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_629
timestamp 1681708930
transform 1 0 1484 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_791
timestamp 1681708930
transform 1 0 1572 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_792
timestamp 1681708930
transform 1 0 1588 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_610
timestamp 1681708930
transform 1 0 1596 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_536
timestamp 1681708930
transform 1 0 1612 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_720
timestamp 1681708930
transform 1 0 1612 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_793
timestamp 1681708930
transform 1 0 1604 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_823
timestamp 1681708930
transform 1 0 1492 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_835
timestamp 1681708930
transform 1 0 1468 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_836
timestamp 1681708930
transform 1 0 1484 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_660
timestamp 1681708930
transform 1 0 1468 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_661
timestamp 1681708930
transform 1 0 1484 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_630
timestamp 1681708930
transform 1 0 1516 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_631
timestamp 1681708930
transform 1 0 1532 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_632
timestamp 1681708930
transform 1 0 1556 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_633
timestamp 1681708930
transform 1 0 1572 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_662
timestamp 1681708930
transform 1 0 1540 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_555
timestamp 1681708930
transform 1 0 1628 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_537
timestamp 1681708930
transform 1 0 1668 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_556
timestamp 1681708930
transform 1 0 1652 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_557
timestamp 1681708930
transform 1 0 1668 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_574
timestamp 1681708930
transform 1 0 1644 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_575
timestamp 1681708930
transform 1 0 1676 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_721
timestamp 1681708930
transform 1 0 1636 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_722
timestamp 1681708930
transform 1 0 1652 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_723
timestamp 1681708930
transform 1 0 1668 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_724
timestamp 1681708930
transform 1 0 1676 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_794
timestamp 1681708930
transform 1 0 1644 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_795
timestamp 1681708930
transform 1 0 1660 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_796
timestamp 1681708930
transform 1 0 1668 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_634
timestamp 1681708930
transform 1 0 1636 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_635
timestamp 1681708930
transform 1 0 1668 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_558
timestamp 1681708930
transform 1 0 1692 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_591
timestamp 1681708930
transform 1 0 1692 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_725
timestamp 1681708930
transform 1 0 1700 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_726
timestamp 1681708930
transform 1 0 1716 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_797
timestamp 1681708930
transform 1 0 1684 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_798
timestamp 1681708930
transform 1 0 1708 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_648
timestamp 1681708930
transform 1 0 1708 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_576
timestamp 1681708930
transform 1 0 1748 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_799
timestamp 1681708930
transform 1 0 1748 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_559
timestamp 1681708930
transform 1 0 1756 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_727
timestamp 1681708930
transform 1 0 1756 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_728
timestamp 1681708930
transform 1 0 1764 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_636
timestamp 1681708930
transform 1 0 1764 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_611
timestamp 1681708930
transform 1 0 1780 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_824
timestamp 1681708930
transform 1 0 1780 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_560
timestamp 1681708930
transform 1 0 1812 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_561
timestamp 1681708930
transform 1 0 1828 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_562
timestamp 1681708930
transform 1 0 1852 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_577
timestamp 1681708930
transform 1 0 1844 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_729
timestamp 1681708930
transform 1 0 1804 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_730
timestamp 1681708930
transform 1 0 1820 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_592
timestamp 1681708930
transform 1 0 1836 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_731
timestamp 1681708930
transform 1 0 1844 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_612
timestamp 1681708930
transform 1 0 1820 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_800
timestamp 1681708930
transform 1 0 1836 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_825
timestamp 1681708930
transform 1 0 1812 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_826
timestamp 1681708930
transform 1 0 1820 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_837
timestamp 1681708930
transform 1 0 1796 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_637
timestamp 1681708930
transform 1 0 1828 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_827
timestamp 1681708930
transform 1 0 1852 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_563
timestamp 1681708930
transform 1 0 1892 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_732
timestamp 1681708930
transform 1 0 1892 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_828
timestamp 1681708930
transform 1 0 1892 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_649
timestamp 1681708930
transform 1 0 1876 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_838
timestamp 1681708930
transform 1 0 1884 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_733
timestamp 1681708930
transform 1 0 1932 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_734
timestamp 1681708930
transform 1 0 1980 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_735
timestamp 1681708930
transform 1 0 1988 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_801
timestamp 1681708930
transform 1 0 1988 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_736
timestamp 1681708930
transform 1 0 2036 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_737
timestamp 1681708930
transform 1 0 2044 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_802
timestamp 1681708930
transform 1 0 2044 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_738
timestamp 1681708930
transform 1 0 2092 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_578
timestamp 1681708930
transform 1 0 2148 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_538
timestamp 1681708930
transform 1 0 2180 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_681
timestamp 1681708930
transform 1 0 2172 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_739
timestamp 1681708930
transform 1 0 2148 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_740
timestamp 1681708930
transform 1 0 2164 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_613
timestamp 1681708930
transform 1 0 2132 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_803
timestamp 1681708930
transform 1 0 2148 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_804
timestamp 1681708930
transform 1 0 2156 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_638
timestamp 1681708930
transform 1 0 2148 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_741
timestamp 1681708930
transform 1 0 2180 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_639
timestamp 1681708930
transform 1 0 2172 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_742
timestamp 1681708930
transform 1 0 2196 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_650
timestamp 1681708930
transform 1 0 2196 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_743
timestamp 1681708930
transform 1 0 2220 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_593
timestamp 1681708930
transform 1 0 2236 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_829
timestamp 1681708930
transform 1 0 2212 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_663
timestamp 1681708930
transform 1 0 2212 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_579
timestamp 1681708930
transform 1 0 2260 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_744
timestamp 1681708930
transform 1 0 2260 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_830
timestamp 1681708930
transform 1 0 2252 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_564
timestamp 1681708930
transform 1 0 2284 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_565
timestamp 1681708930
transform 1 0 2332 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_580
timestamp 1681708930
transform 1 0 2340 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_594
timestamp 1681708930
transform 1 0 2308 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_595
timestamp 1681708930
transform 1 0 2324 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_745
timestamp 1681708930
transform 1 0 2332 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_805
timestamp 1681708930
transform 1 0 2284 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_614
timestamp 1681708930
transform 1 0 2292 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_806
timestamp 1681708930
transform 1 0 2308 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_807
timestamp 1681708930
transform 1 0 2332 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_831
timestamp 1681708930
transform 1 0 2292 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_672
timestamp 1681708930
transform 1 0 2284 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_832
timestamp 1681708930
transform 1 0 2324 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_839
timestamp 1681708930
transform 1 0 2308 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_840
timestamp 1681708930
transform 1 0 2316 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_651
timestamp 1681708930
transform 1 0 2324 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_664
timestamp 1681708930
transform 1 0 2316 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_746
timestamp 1681708930
transform 1 0 2356 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_808
timestamp 1681708930
transform 1 0 2348 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_615
timestamp 1681708930
transform 1 0 2356 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_596
timestamp 1681708930
transform 1 0 2380 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_566
timestamp 1681708930
transform 1 0 2412 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_682
timestamp 1681708930
transform 1 0 2404 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_683
timestamp 1681708930
transform 1 0 2412 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_747
timestamp 1681708930
transform 1 0 2388 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_748
timestamp 1681708930
transform 1 0 2396 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_749
timestamp 1681708930
transform 1 0 2412 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_809
timestamp 1681708930
transform 1 0 2380 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_616
timestamp 1681708930
transform 1 0 2388 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_617
timestamp 1681708930
transform 1 0 2412 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_833
timestamp 1681708930
transform 1 0 2380 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_652
timestamp 1681708930
transform 1 0 2380 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_653
timestamp 1681708930
transform 1 0 2404 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_567
timestamp 1681708930
transform 1 0 2484 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_539
timestamp 1681708930
transform 1 0 2516 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_581
timestamp 1681708930
transform 1 0 2500 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_750
timestamp 1681708930
transform 1 0 2492 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_751
timestamp 1681708930
transform 1 0 2500 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_810
timestamp 1681708930
transform 1 0 2468 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_811
timestamp 1681708930
transform 1 0 2500 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_640
timestamp 1681708930
transform 1 0 2468 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_540
timestamp 1681708930
transform 1 0 2612 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_568
timestamp 1681708930
transform 1 0 2596 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_752
timestamp 1681708930
transform 1 0 2548 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_753
timestamp 1681708930
transform 1 0 2556 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_812
timestamp 1681708930
transform 1 0 2548 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_678
timestamp 1681708930
transform 1 0 2668 0 1 2155
box -2 -2 2 2
use M2_M1  M2_M1_754
timestamp 1681708930
transform 1 0 2604 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_597
timestamp 1681708930
transform 1 0 2660 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_755
timestamp 1681708930
transform 1 0 2732 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_813
timestamp 1681708930
transform 1 0 2604 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_814
timestamp 1681708930
transform 1 0 2636 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_641
timestamp 1681708930
transform 1 0 2604 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_642
timestamp 1681708930
transform 1 0 2668 0 1 2115
box -3 -3 3 3
use top_mod_new_VIA0  top_mod_new_VIA0_10
timestamp 1681708930
transform 1 0 24 0 1 2070
box -10 -3 10 3
use INVX2  INVX2_38
timestamp 1681708930
transform 1 0 72 0 -1 2170
box -9 -3 26 105
use FILL  FILL_185
timestamp 1681708930
transform 1 0 88 0 -1 2170
box -8 -3 16 105
use FILL  FILL_186
timestamp 1681708930
transform 1 0 96 0 -1 2170
box -8 -3 16 105
use FILL  FILL_187
timestamp 1681708930
transform 1 0 104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_188
timestamp 1681708930
transform 1 0 112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_189
timestamp 1681708930
transform 1 0 120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_190
timestamp 1681708930
transform 1 0 128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_191
timestamp 1681708930
transform 1 0 136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_192
timestamp 1681708930
transform 1 0 144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_193
timestamp 1681708930
transform 1 0 152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_194
timestamp 1681708930
transform 1 0 160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_195
timestamp 1681708930
transform 1 0 168 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_9
timestamp 1681708930
transform -1 0 216 0 -1 2170
box -8 -3 46 105
use FILL  FILL_196
timestamp 1681708930
transform 1 0 216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_197
timestamp 1681708930
transform 1 0 224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_198
timestamp 1681708930
transform 1 0 232 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_42
timestamp 1681708930
transform -1 0 256 0 -1 2170
box -9 -3 26 105
use OAI22X1  OAI22X1_10
timestamp 1681708930
transform -1 0 296 0 -1 2170
box -8 -3 46 105
use FILL  FILL_199
timestamp 1681708930
transform 1 0 296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_201
timestamp 1681708930
transform 1 0 304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_203
timestamp 1681708930
transform 1 0 312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_210
timestamp 1681708930
transform 1 0 320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_211
timestamp 1681708930
transform 1 0 328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_212
timestamp 1681708930
transform 1 0 336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_213
timestamp 1681708930
transform 1 0 344 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_16
timestamp 1681708930
transform 1 0 352 0 -1 2170
box -8 -3 104 105
use FILL  FILL_214
timestamp 1681708930
transform 1 0 448 0 -1 2170
box -8 -3 16 105
use FILL  FILL_233
timestamp 1681708930
transform 1 0 456 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_49
timestamp 1681708930
transform 1 0 464 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_50
timestamp 1681708930
transform 1 0 480 0 -1 2170
box -9 -3 26 105
use FILL  FILL_234
timestamp 1681708930
transform 1 0 496 0 -1 2170
box -8 -3 16 105
use FILL  FILL_235
timestamp 1681708930
transform 1 0 504 0 -1 2170
box -8 -3 16 105
use FILL  FILL_236
timestamp 1681708930
transform 1 0 512 0 -1 2170
box -8 -3 16 105
use FILL  FILL_237
timestamp 1681708930
transform 1 0 520 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_673
timestamp 1681708930
transform 1 0 572 0 1 2075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_17
timestamp 1681708930
transform 1 0 528 0 -1 2170
box -8 -3 104 105
use M3_M2  M3_M2_674
timestamp 1681708930
transform 1 0 652 0 1 2075
box -3 -3 3 3
use XOR2X1  XOR2X1_16
timestamp 1681708930
transform -1 0 680 0 -1 2170
box -8 -3 64 105
use NAND3X1  NAND3X1_19
timestamp 1681708930
transform 1 0 680 0 -1 2170
box -8 -3 40 105
use XOR2X1  XOR2X1_17
timestamp 1681708930
transform -1 0 768 0 -1 2170
box -8 -3 64 105
use FILL  FILL_238
timestamp 1681708930
transform 1 0 768 0 -1 2170
box -8 -3 16 105
use FILL  FILL_239
timestamp 1681708930
transform 1 0 776 0 -1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_20
timestamp 1681708930
transform 1 0 784 0 -1 2170
box -8 -3 34 105
use FILL  FILL_240
timestamp 1681708930
transform 1 0 816 0 -1 2170
box -8 -3 16 105
use FILL  FILL_241
timestamp 1681708930
transform 1 0 824 0 -1 2170
box -8 -3 16 105
use FILL  FILL_242
timestamp 1681708930
transform 1 0 832 0 -1 2170
box -8 -3 16 105
use FILL  FILL_243
timestamp 1681708930
transform 1 0 840 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_21
timestamp 1681708930
transform 1 0 848 0 -1 2170
box -8 -3 104 105
use FILL  FILL_272
timestamp 1681708930
transform 1 0 944 0 -1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_21
timestamp 1681708930
transform 1 0 952 0 -1 2170
box -8 -3 32 105
use FILL  FILL_273
timestamp 1681708930
transform 1 0 976 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_22
timestamp 1681708930
transform 1 0 984 0 -1 2170
box -8 -3 104 105
use OAI21X1  OAI21X1_25
timestamp 1681708930
transform -1 0 1112 0 -1 2170
box -8 -3 34 105
use XOR2X1  XOR2X1_19
timestamp 1681708930
transform -1 0 1168 0 -1 2170
box -8 -3 64 105
use NAND2X1  NAND2X1_22
timestamp 1681708930
transform 1 0 1168 0 -1 2170
box -8 -3 32 105
use FILL  FILL_274
timestamp 1681708930
transform 1 0 1192 0 -1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_26
timestamp 1681708930
transform 1 0 1200 0 -1 2170
box -8 -3 34 105
use FILL  FILL_275
timestamp 1681708930
transform 1 0 1232 0 -1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_23
timestamp 1681708930
transform -1 0 1264 0 -1 2170
box -8 -3 32 105
use FILL  FILL_276
timestamp 1681708930
transform 1 0 1264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_277
timestamp 1681708930
transform 1 0 1272 0 -1 2170
box -8 -3 16 105
use XOR2X1  XOR2X1_20
timestamp 1681708930
transform -1 0 1336 0 -1 2170
box -8 -3 64 105
use M3_M2  M3_M2_675
timestamp 1681708930
transform 1 0 1364 0 1 2075
box -3 -3 3 3
use XOR2X1  XOR2X1_21
timestamp 1681708930
transform -1 0 1392 0 -1 2170
box -8 -3 64 105
use XOR2X1  XOR2X1_22
timestamp 1681708930
transform -1 0 1448 0 -1 2170
box -8 -3 64 105
use INVX2  INVX2_54
timestamp 1681708930
transform -1 0 1464 0 -1 2170
box -9 -3 26 105
use NAND3X1  NAND3X1_22
timestamp 1681708930
transform 1 0 1464 0 -1 2170
box -8 -3 40 105
use AOI22X1  AOI22X1_5
timestamp 1681708930
transform 1 0 1496 0 -1 2170
box -8 -3 46 105
use OR2X1  OR2X1_4
timestamp 1681708930
transform -1 0 1568 0 -1 2170
box -8 -3 40 105
use AOI22X1  AOI22X1_6
timestamp 1681708930
transform -1 0 1608 0 -1 2170
box -8 -3 46 105
use FILL  FILL_278
timestamp 1681708930
transform 1 0 1608 0 -1 2170
box -8 -3 16 105
use FILL  FILL_279
timestamp 1681708930
transform 1 0 1616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_280
timestamp 1681708930
transform 1 0 1624 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_13
timestamp 1681708930
transform -1 0 1672 0 -1 2170
box -8 -3 46 105
use FILL  FILL_281
timestamp 1681708930
transform 1 0 1672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_282
timestamp 1681708930
transform 1 0 1680 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_7
timestamp 1681708930
transform 1 0 1688 0 -1 2170
box -8 -3 46 105
use INVX2  INVX2_55
timestamp 1681708930
transform -1 0 1744 0 -1 2170
box -9 -3 26 105
use FILL  FILL_283
timestamp 1681708930
transform 1 0 1744 0 -1 2170
box -8 -3 16 105
use FILL  FILL_284
timestamp 1681708930
transform 1 0 1752 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_56
timestamp 1681708930
transform 1 0 1760 0 -1 2170
box -9 -3 26 105
use FILL  FILL_285
timestamp 1681708930
transform 1 0 1776 0 -1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_23
timestamp 1681708930
transform -1 0 1816 0 -1 2170
box -8 -3 40 105
use OAI21X1  OAI21X1_27
timestamp 1681708930
transform -1 0 1848 0 -1 2170
box -8 -3 34 105
use FILL  FILL_286
timestamp 1681708930
transform 1 0 1848 0 -1 2170
box -8 -3 16 105
use FILL  FILL_296
timestamp 1681708930
transform 1 0 1856 0 -1 2170
box -8 -3 16 105
use FILL  FILL_297
timestamp 1681708930
transform 1 0 1864 0 -1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_25
timestamp 1681708930
transform -1 0 1904 0 -1 2170
box -8 -3 40 105
use FILL  FILL_298
timestamp 1681708930
transform 1 0 1904 0 -1 2170
box -8 -3 16 105
use FILL  FILL_299
timestamp 1681708930
transform 1 0 1912 0 -1 2170
box -8 -3 16 105
use FILL  FILL_300
timestamp 1681708930
transform 1 0 1920 0 -1 2170
box -8 -3 16 105
use XOR2X1  XOR2X1_27
timestamp 1681708930
transform 1 0 1928 0 -1 2170
box -8 -3 64 105
use XOR2X1  XOR2X1_28
timestamp 1681708930
transform 1 0 1984 0 -1 2170
box -8 -3 64 105
use XOR2X1  XOR2X1_29
timestamp 1681708930
transform 1 0 2040 0 -1 2170
box -8 -3 64 105
use XOR2X1  XOR2X1_30
timestamp 1681708930
transform 1 0 2096 0 -1 2170
box -8 -3 64 105
use NOR2X1  NOR2X1_17
timestamp 1681708930
transform -1 0 2176 0 -1 2170
box -8 -3 32 105
use M3_M2  M3_M2_676
timestamp 1681708930
transform 1 0 2188 0 1 2075
box -3 -3 3 3
use FILL  FILL_301
timestamp 1681708930
transform 1 0 2176 0 -1 2170
box -8 -3 16 105
use FILL  FILL_303
timestamp 1681708930
transform 1 0 2184 0 -1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_26
timestamp 1681708930
transform 1 0 2192 0 -1 2170
box -8 -3 32 105
use OAI21X1  OAI21X1_28
timestamp 1681708930
transform 1 0 2216 0 -1 2170
box -8 -3 34 105
use FILL  FILL_305
timestamp 1681708930
transform 1 0 2248 0 -1 2170
box -8 -3 16 105
use FILL  FILL_306
timestamp 1681708930
transform 1 0 2256 0 -1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_26
timestamp 1681708930
transform -1 0 2296 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_27
timestamp 1681708930
transform 1 0 2296 0 -1 2170
box -8 -3 40 105
use INVX2  INVX2_58
timestamp 1681708930
transform 1 0 2328 0 -1 2170
box -9 -3 26 105
use FILL  FILL_307
timestamp 1681708930
transform 1 0 2344 0 -1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_30
timestamp 1681708930
transform 1 0 2352 0 -1 2170
box -8 -3 34 105
use NOR2X1  NOR2X1_18
timestamp 1681708930
transform -1 0 2408 0 -1 2170
box -8 -3 32 105
use OR2X1  OR2X1_5
timestamp 1681708930
transform 1 0 2408 0 -1 2170
box -8 -3 40 105
use XOR2X1  XOR2X1_33
timestamp 1681708930
transform -1 0 2496 0 -1 2170
box -8 -3 64 105
use XOR2X1  XOR2X1_34
timestamp 1681708930
transform -1 0 2552 0 -1 2170
box -8 -3 64 105
use XOR2X1  XOR2X1_35
timestamp 1681708930
transform -1 0 2608 0 -1 2170
box -8 -3 64 105
use XOR2X1  XOR2X1_36
timestamp 1681708930
transform 1 0 2608 0 -1 2170
box -8 -3 64 105
use top_mod_new_VIA0  top_mod_new_VIA0_11
timestamp 1681708930
transform 1 0 2712 0 1 2070
box -10 -3 10 3
use M2_M1  M2_M1_857
timestamp 1681708930
transform 1 0 76 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_858
timestamp 1681708930
transform 1 0 140 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_920
timestamp 1681708930
transform 1 0 164 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_859
timestamp 1681708930
transform 1 0 212 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_860
timestamp 1681708930
transform 1 0 236 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_921
timestamp 1681708930
transform 1 0 212 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_922
timestamp 1681708930
transform 1 0 228 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_923
timestamp 1681708930
transform 1 0 244 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_793
timestamp 1681708930
transform 1 0 212 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_781
timestamp 1681708930
transform 1 0 244 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_694
timestamp 1681708930
transform 1 0 276 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_695
timestamp 1681708930
transform 1 0 364 0 1 2045
box -3 -3 3 3
use M2_M1  M2_M1_861
timestamp 1681708930
transform 1 0 300 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_862
timestamp 1681708930
transform 1 0 356 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_863
timestamp 1681708930
transform 1 0 372 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_864
timestamp 1681708930
transform 1 0 388 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_924
timestamp 1681708930
transform 1 0 276 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_925
timestamp 1681708930
transform 1 0 364 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_926
timestamp 1681708930
transform 1 0 380 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_782
timestamp 1681708930
transform 1 0 340 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_783
timestamp 1681708930
transform 1 0 356 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_784
timestamp 1681708930
transform 1 0 372 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_794
timestamp 1681708930
transform 1 0 268 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_785
timestamp 1681708930
transform 1 0 412 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_706
timestamp 1681708930
transform 1 0 428 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_927
timestamp 1681708930
transform 1 0 428 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_928
timestamp 1681708930
transform 1 0 436 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_764
timestamp 1681708930
transform 1 0 444 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_991
timestamp 1681708930
transform 1 0 444 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_795
timestamp 1681708930
transform 1 0 452 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_865
timestamp 1681708930
transform 1 0 468 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_866
timestamp 1681708930
transform 1 0 484 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_765
timestamp 1681708930
transform 1 0 468 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_929
timestamp 1681708930
transform 1 0 476 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_766
timestamp 1681708930
transform 1 0 484 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_930
timestamp 1681708930
transform 1 0 500 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_685
timestamp 1681708930
transform 1 0 564 0 1 2055
box -3 -3 3 3
use M2_M1  M2_M1_867
timestamp 1681708930
transform 1 0 540 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_868
timestamp 1681708930
transform 1 0 596 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_869
timestamp 1681708930
transform 1 0 604 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_931
timestamp 1681708930
transform 1 0 516 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_767
timestamp 1681708930
transform 1 0 540 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_768
timestamp 1681708930
transform 1 0 596 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_786
timestamp 1681708930
transform 1 0 516 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_787
timestamp 1681708930
transform 1 0 580 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_796
timestamp 1681708930
transform 1 0 516 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_696
timestamp 1681708930
transform 1 0 628 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_752
timestamp 1681708930
transform 1 0 620 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_932
timestamp 1681708930
transform 1 0 620 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_707
timestamp 1681708930
transform 1 0 636 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_844
timestamp 1681708930
transform 1 0 644 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_841
timestamp 1681708930
transform 1 0 676 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_845
timestamp 1681708930
transform 1 0 692 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_753
timestamp 1681708930
transform 1 0 676 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_870
timestamp 1681708930
transform 1 0 684 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_871
timestamp 1681708930
transform 1 0 700 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_769
timestamp 1681708930
transform 1 0 692 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_933
timestamp 1681708930
transform 1 0 700 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_788
timestamp 1681708930
transform 1 0 684 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_727
timestamp 1681708930
transform 1 0 740 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_677
timestamp 1681708930
transform 1 0 764 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_678
timestamp 1681708930
transform 1 0 788 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_708
timestamp 1681708930
transform 1 0 780 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_754
timestamp 1681708930
transform 1 0 772 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_728
timestamp 1681708930
transform 1 0 788 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_686
timestamp 1681708930
transform 1 0 1012 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_697
timestamp 1681708930
transform 1 0 996 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_709
timestamp 1681708930
transform 1 0 892 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_710
timestamp 1681708930
transform 1 0 972 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_846
timestamp 1681708930
transform 1 0 796 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1681708930
transform 1 0 788 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_934
timestamp 1681708930
transform 1 0 772 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_935
timestamp 1681708930
transform 1 0 780 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_729
timestamp 1681708930
transform 1 0 812 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_847
timestamp 1681708930
transform 1 0 996 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_873
timestamp 1681708930
transform 1 0 836 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_874
timestamp 1681708930
transform 1 0 892 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_875
timestamp 1681708930
transform 1 0 956 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_755
timestamp 1681708930
transform 1 0 980 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_876
timestamp 1681708930
transform 1 0 988 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_770
timestamp 1681708930
transform 1 0 796 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_936
timestamp 1681708930
transform 1 0 812 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_771
timestamp 1681708930
transform 1 0 860 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_772
timestamp 1681708930
transform 1 0 892 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_937
timestamp 1681708930
transform 1 0 908 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_938
timestamp 1681708930
transform 1 0 996 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_789
timestamp 1681708930
transform 1 0 796 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_797
timestamp 1681708930
transform 1 0 812 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_798
timestamp 1681708930
transform 1 0 852 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_799
timestamp 1681708930
transform 1 0 876 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_790
timestamp 1681708930
transform 1 0 956 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_791
timestamp 1681708930
transform 1 0 996 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_800
timestamp 1681708930
transform 1 0 908 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_801
timestamp 1681708930
transform 1 0 980 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_679
timestamp 1681708930
transform 1 0 1092 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_877
timestamp 1681708930
transform 1 0 1028 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_878
timestamp 1681708930
transform 1 0 1044 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_939
timestamp 1681708930
transform 1 0 1020 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_940
timestamp 1681708930
transform 1 0 1028 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_756
timestamp 1681708930
transform 1 0 1076 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_879
timestamp 1681708930
transform 1 0 1084 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_941
timestamp 1681708930
transform 1 0 1076 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_687
timestamp 1681708930
transform 1 0 1116 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_711
timestamp 1681708930
transform 1 0 1100 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_848
timestamp 1681708930
transform 1 0 1100 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_730
timestamp 1681708930
transform 1 0 1108 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_942
timestamp 1681708930
transform 1 0 1100 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_680
timestamp 1681708930
transform 1 0 1220 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_698
timestamp 1681708930
transform 1 0 1188 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_712
timestamp 1681708930
transform 1 0 1180 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_731
timestamp 1681708930
transform 1 0 1188 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_757
timestamp 1681708930
transform 1 0 1156 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_880
timestamp 1681708930
transform 1 0 1180 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_881
timestamp 1681708930
transform 1 0 1188 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_943
timestamp 1681708930
transform 1 0 1156 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_944
timestamp 1681708930
transform 1 0 1164 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_688
timestamp 1681708930
transform 1 0 1260 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_699
timestamp 1681708930
transform 1 0 1300 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_713
timestamp 1681708930
transform 1 0 1300 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_689
timestamp 1681708930
transform 1 0 1340 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_714
timestamp 1681708930
transform 1 0 1340 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_732
timestamp 1681708930
transform 1 0 1308 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_681
timestamp 1681708930
transform 1 0 1420 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_715
timestamp 1681708930
transform 1 0 1396 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_733
timestamp 1681708930
transform 1 0 1364 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_882
timestamp 1681708930
transform 1 0 1252 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_883
timestamp 1681708930
transform 1 0 1308 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_884
timestamp 1681708930
transform 1 0 1340 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_945
timestamp 1681708930
transform 1 0 1212 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_946
timestamp 1681708930
transform 1 0 1228 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_802
timestamp 1681708930
transform 1 0 1212 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_773
timestamp 1681708930
transform 1 0 1308 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_947
timestamp 1681708930
transform 1 0 1316 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_690
timestamp 1681708930
transform 1 0 1444 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_700
timestamp 1681708930
transform 1 0 1452 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_691
timestamp 1681708930
transform 1 0 1492 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_692
timestamp 1681708930
transform 1 0 1524 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_716
timestamp 1681708930
transform 1 0 1476 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_717
timestamp 1681708930
transform 1 0 1492 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_842
timestamp 1681708930
transform 1 0 1500 0 1 2035
box -2 -2 2 2
use M3_M2  M3_M2_718
timestamp 1681708930
transform 1 0 1516 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_734
timestamp 1681708930
transform 1 0 1428 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_735
timestamp 1681708930
transform 1 0 1444 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_736
timestamp 1681708930
transform 1 0 1460 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_758
timestamp 1681708930
transform 1 0 1396 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_885
timestamp 1681708930
transform 1 0 1420 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_886
timestamp 1681708930
transform 1 0 1460 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_948
timestamp 1681708930
transform 1 0 1364 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_949
timestamp 1681708930
transform 1 0 1372 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_803
timestamp 1681708930
transform 1 0 1308 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_804
timestamp 1681708930
transform 1 0 1356 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_950
timestamp 1681708930
transform 1 0 1420 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_951
timestamp 1681708930
transform 1 0 1428 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_849
timestamp 1681708930
transform 1 0 1492 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_737
timestamp 1681708930
transform 1 0 1500 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_850
timestamp 1681708930
transform 1 0 1508 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_851
timestamp 1681708930
transform 1 0 1516 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_887
timestamp 1681708930
transform 1 0 1492 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_952
timestamp 1681708930
transform 1 0 1476 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_843
timestamp 1681708930
transform 1 0 1540 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_852
timestamp 1681708930
transform 1 0 1540 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_888
timestamp 1681708930
transform 1 0 1532 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_774
timestamp 1681708930
transform 1 0 1516 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_775
timestamp 1681708930
transform 1 0 1540 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_953
timestamp 1681708930
transform 1 0 1548 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_693
timestamp 1681708930
transform 1 0 1564 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_701
timestamp 1681708930
transform 1 0 1564 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_719
timestamp 1681708930
transform 1 0 1588 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_738
timestamp 1681708930
transform 1 0 1580 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_720
timestamp 1681708930
transform 1 0 1612 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_889
timestamp 1681708930
transform 1 0 1556 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_890
timestamp 1681708930
transform 1 0 1564 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_891
timestamp 1681708930
transform 1 0 1580 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_892
timestamp 1681708930
transform 1 0 1596 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_893
timestamp 1681708930
transform 1 0 1604 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_954
timestamp 1681708930
transform 1 0 1572 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_955
timestamp 1681708930
transform 1 0 1588 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_805
timestamp 1681708930
transform 1 0 1572 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_721
timestamp 1681708930
transform 1 0 1652 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_894
timestamp 1681708930
transform 1 0 1636 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_759
timestamp 1681708930
transform 1 0 1644 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_776
timestamp 1681708930
transform 1 0 1620 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_956
timestamp 1681708930
transform 1 0 1628 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_777
timestamp 1681708930
transform 1 0 1636 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_957
timestamp 1681708930
transform 1 0 1644 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_992
timestamp 1681708930
transform 1 0 1620 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_806
timestamp 1681708930
transform 1 0 1628 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_958
timestamp 1681708930
transform 1 0 1692 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_722
timestamp 1681708930
transform 1 0 1708 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_993
timestamp 1681708930
transform 1 0 1700 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_959
timestamp 1681708930
transform 1 0 1724 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_807
timestamp 1681708930
transform 1 0 1724 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_960
timestamp 1681708930
transform 1 0 1740 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_723
timestamp 1681708930
transform 1 0 1780 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_853
timestamp 1681708930
transform 1 0 1780 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_682
timestamp 1681708930
transform 1 0 1796 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_895
timestamp 1681708930
transform 1 0 1788 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_760
timestamp 1681708930
transform 1 0 1796 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_896
timestamp 1681708930
transform 1 0 1820 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_961
timestamp 1681708930
transform 1 0 1796 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_962
timestamp 1681708930
transform 1 0 1804 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_963
timestamp 1681708930
transform 1 0 1812 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_778
timestamp 1681708930
transform 1 0 1820 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_964
timestamp 1681708930
transform 1 0 1828 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_808
timestamp 1681708930
transform 1 0 1804 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_683
timestamp 1681708930
transform 1 0 1876 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_761
timestamp 1681708930
transform 1 0 1868 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_965
timestamp 1681708930
transform 1 0 1868 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_739
timestamp 1681708930
transform 1 0 1884 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_684
timestamp 1681708930
transform 1 0 1908 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_724
timestamp 1681708930
transform 1 0 1916 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_740
timestamp 1681708930
transform 1 0 1924 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_897
timestamp 1681708930
transform 1 0 1884 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_898
timestamp 1681708930
transform 1 0 1892 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_899
timestamp 1681708930
transform 1 0 1908 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_900
timestamp 1681708930
transform 1 0 1924 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_779
timestamp 1681708930
transform 1 0 1892 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_966
timestamp 1681708930
transform 1 0 1916 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_967
timestamp 1681708930
transform 1 0 1940 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_809
timestamp 1681708930
transform 1 0 1980 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_741
timestamp 1681708930
transform 1 0 2012 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_901
timestamp 1681708930
transform 1 0 2012 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1681708930
transform 1 0 2060 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_968
timestamp 1681708930
transform 1 0 2036 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_969
timestamp 1681708930
transform 1 0 2052 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_994
timestamp 1681708930
transform 1 0 2060 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_810
timestamp 1681708930
transform 1 0 2028 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_742
timestamp 1681708930
transform 1 0 2076 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_903
timestamp 1681708930
transform 1 0 2076 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_970
timestamp 1681708930
transform 1 0 2108 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_702
timestamp 1681708930
transform 1 0 2124 0 1 2045
box -3 -3 3 3
use M2_M1  M2_M1_904
timestamp 1681708930
transform 1 0 2124 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_971
timestamp 1681708930
transform 1 0 2116 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_743
timestamp 1681708930
transform 1 0 2156 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_972
timestamp 1681708930
transform 1 0 2148 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_703
timestamp 1681708930
transform 1 0 2164 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_744
timestamp 1681708930
transform 1 0 2188 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_745
timestamp 1681708930
transform 1 0 2228 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_905
timestamp 1681708930
transform 1 0 2188 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_973
timestamp 1681708930
transform 1 0 2172 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_995
timestamp 1681708930
transform 1 0 2164 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_811
timestamp 1681708930
transform 1 0 2164 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_906
timestamp 1681708930
transform 1 0 2236 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_907
timestamp 1681708930
transform 1 0 2252 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_974
timestamp 1681708930
transform 1 0 2220 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_975
timestamp 1681708930
transform 1 0 2228 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_976
timestamp 1681708930
transform 1 0 2252 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_812
timestamp 1681708930
transform 1 0 2252 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_854
timestamp 1681708930
transform 1 0 2260 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_746
timestamp 1681708930
transform 1 0 2300 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_908
timestamp 1681708930
transform 1 0 2292 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_909
timestamp 1681708930
transform 1 0 2300 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_977
timestamp 1681708930
transform 1 0 2284 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_747
timestamp 1681708930
transform 1 0 2324 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_978
timestamp 1681708930
transform 1 0 2308 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_910
timestamp 1681708930
transform 1 0 2324 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_996
timestamp 1681708930
transform 1 0 2324 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_813
timestamp 1681708930
transform 1 0 2324 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_725
timestamp 1681708930
transform 1 0 2364 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_748
timestamp 1681708930
transform 1 0 2380 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_911
timestamp 1681708930
transform 1 0 2348 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_912
timestamp 1681708930
transform 1 0 2372 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_979
timestamp 1681708930
transform 1 0 2340 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_980
timestamp 1681708930
transform 1 0 2356 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_981
timestamp 1681708930
transform 1 0 2372 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_982
timestamp 1681708930
transform 1 0 2388 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_814
timestamp 1681708930
transform 1 0 2356 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_704
timestamp 1681708930
transform 1 0 2436 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_726
timestamp 1681708930
transform 1 0 2444 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_855
timestamp 1681708930
transform 1 0 2444 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_913
timestamp 1681708930
transform 1 0 2444 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_983
timestamp 1681708930
transform 1 0 2436 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_749
timestamp 1681708930
transform 1 0 2468 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_984
timestamp 1681708930
transform 1 0 2460 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_985
timestamp 1681708930
transform 1 0 2468 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_856
timestamp 1681708930
transform 1 0 2492 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_750
timestamp 1681708930
transform 1 0 2532 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_705
timestamp 1681708930
transform 1 0 2580 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_751
timestamp 1681708930
transform 1 0 2644 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_914
timestamp 1681708930
transform 1 0 2532 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_915
timestamp 1681708930
transform 1 0 2548 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_916
timestamp 1681708930
transform 1 0 2580 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_917
timestamp 1681708930
transform 1 0 2604 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_986
timestamp 1681708930
transform 1 0 2492 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_987
timestamp 1681708930
transform 1 0 2500 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_988
timestamp 1681708930
transform 1 0 2548 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_792
timestamp 1681708930
transform 1 0 2500 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_815
timestamp 1681708930
transform 1 0 2532 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_762
timestamp 1681708930
transform 1 0 2612 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_763
timestamp 1681708930
transform 1 0 2636 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_918
timestamp 1681708930
transform 1 0 2644 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_919
timestamp 1681708930
transform 1 0 2660 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_989
timestamp 1681708930
transform 1 0 2604 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_780
timestamp 1681708930
transform 1 0 2660 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_990
timestamp 1681708930
transform 1 0 2668 0 1 2005
box -2 -2 2 2
use top_mod_new_VIA0  top_mod_new_VIA0_12
timestamp 1681708930
transform 1 0 48 0 1 1970
box -10 -3 10 3
use FILL  FILL_313
timestamp 1681708930
transform 1 0 72 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_816
timestamp 1681708930
transform 1 0 164 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_23
timestamp 1681708930
transform -1 0 176 0 1 1970
box -8 -3 104 105
use FILL  FILL_314
timestamp 1681708930
transform 1 0 176 0 1 1970
box -8 -3 16 105
use FILL  FILL_315
timestamp 1681708930
transform 1 0 184 0 1 1970
box -8 -3 16 105
use FILL  FILL_316
timestamp 1681708930
transform 1 0 192 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_817
timestamp 1681708930
transform 1 0 212 0 1 1975
box -3 -3 3 3
use FILL  FILL_317
timestamp 1681708930
transform 1 0 200 0 1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_14
timestamp 1681708930
transform 1 0 208 0 1 1970
box -8 -3 46 105
use FILL  FILL_318
timestamp 1681708930
transform 1 0 248 0 1 1970
box -8 -3 16 105
use FILL  FILL_319
timestamp 1681708930
transform 1 0 256 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_818
timestamp 1681708930
transform 1 0 276 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_24
timestamp 1681708930
transform 1 0 264 0 1 1970
box -8 -3 104 105
use M3_M2  M3_M2_819
timestamp 1681708930
transform 1 0 372 0 1 1975
box -3 -3 3 3
use OAI22X1  OAI22X1_15
timestamp 1681708930
transform -1 0 400 0 1 1970
box -8 -3 46 105
use FILL  FILL_320
timestamp 1681708930
transform 1 0 400 0 1 1970
box -8 -3 16 105
use FILL  FILL_321
timestamp 1681708930
transform 1 0 408 0 1 1970
box -8 -3 16 105
use FILL  FILL_322
timestamp 1681708930
transform 1 0 416 0 1 1970
box -8 -3 16 105
use FILL  FILL_323
timestamp 1681708930
transform 1 0 424 0 1 1970
box -8 -3 16 105
use FILL  FILL_324
timestamp 1681708930
transform 1 0 432 0 1 1970
box -8 -3 16 105
use FILL  FILL_325
timestamp 1681708930
transform 1 0 440 0 1 1970
box -8 -3 16 105
use FILL  FILL_326
timestamp 1681708930
transform 1 0 448 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_820
timestamp 1681708930
transform 1 0 492 0 1 1975
box -3 -3 3 3
use OAI22X1  OAI22X1_16
timestamp 1681708930
transform -1 0 496 0 1 1970
box -8 -3 46 105
use M3_M2  M3_M2_821
timestamp 1681708930
transform 1 0 508 0 1 1975
box -3 -3 3 3
use FILL  FILL_327
timestamp 1681708930
transform 1 0 496 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_25
timestamp 1681708930
transform 1 0 504 0 1 1970
box -8 -3 104 105
use M3_M2  M3_M2_822
timestamp 1681708930
transform 1 0 612 0 1 1975
box -3 -3 3 3
use FILL  FILL_328
timestamp 1681708930
transform 1 0 600 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_61
timestamp 1681708930
transform -1 0 624 0 1 1970
box -9 -3 26 105
use FILL  FILL_329
timestamp 1681708930
transform 1 0 624 0 1 1970
box -8 -3 16 105
use FILL  FILL_330
timestamp 1681708930
transform 1 0 632 0 1 1970
box -8 -3 16 105
use FILL  FILL_331
timestamp 1681708930
transform 1 0 640 0 1 1970
box -8 -3 16 105
use FILL  FILL_335
timestamp 1681708930
transform 1 0 648 0 1 1970
box -8 -3 16 105
use FILL  FILL_337
timestamp 1681708930
transform 1 0 656 0 1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_30
timestamp 1681708930
transform -1 0 696 0 1 1970
box -8 -3 40 105
use M3_M2  M3_M2_823
timestamp 1681708930
transform 1 0 708 0 1 1975
box -3 -3 3 3
use FILL  FILL_338
timestamp 1681708930
transform 1 0 696 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_824
timestamp 1681708930
transform 1 0 756 0 1 1975
box -3 -3 3 3
use XOR2X1  XOR2X1_37
timestamp 1681708930
transform -1 0 760 0 1 1970
box -8 -3 64 105
use FILL  FILL_339
timestamp 1681708930
transform 1 0 760 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_825
timestamp 1681708930
transform 1 0 780 0 1 1975
box -3 -3 3 3
use FILL  FILL_340
timestamp 1681708930
transform 1 0 768 0 1 1970
box -8 -3 16 105
use NAND2X1  NAND2X1_28
timestamp 1681708930
transform 1 0 776 0 1 1970
box -8 -3 32 105
use M3_M2  M3_M2_826
timestamp 1681708930
transform 1 0 820 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_827
timestamp 1681708930
transform 1 0 884 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_28
timestamp 1681708930
transform 1 0 800 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_29
timestamp 1681708930
transform 1 0 896 0 1 1970
box -8 -3 104 105
use OAI21X1  OAI21X1_33
timestamp 1681708930
transform -1 0 1024 0 1 1970
box -8 -3 34 105
use XOR2X1  XOR2X1_38
timestamp 1681708930
transform -1 0 1080 0 1 1970
box -8 -3 64 105
use NAND2X1  NAND2X1_29
timestamp 1681708930
transform 1 0 1080 0 1 1970
box -8 -3 32 105
use XOR2X1  XOR2X1_39
timestamp 1681708930
transform 1 0 1104 0 1 1970
box -8 -3 64 105
use XOR2X1  XOR2X1_40
timestamp 1681708930
transform -1 0 1216 0 1 1970
box -8 -3 64 105
use DFFNEGX1  DFFNEGX1_30
timestamp 1681708930
transform 1 0 1216 0 1 1970
box -8 -3 104 105
use XOR2X1  XOR2X1_41
timestamp 1681708930
transform -1 0 1368 0 1 1970
box -8 -3 64 105
use XOR2X1  XOR2X1_42
timestamp 1681708930
transform 1 0 1368 0 1 1970
box -8 -3 64 105
use XOR2X1  XOR2X1_43
timestamp 1681708930
transform 1 0 1424 0 1 1970
box -8 -3 64 105
use NAND3X1  NAND3X1_31
timestamp 1681708930
transform 1 0 1480 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_32
timestamp 1681708930
transform -1 0 1544 0 1 1970
box -8 -3 40 105
use INVX2  INVX2_66
timestamp 1681708930
transform 1 0 1544 0 1 1970
box -9 -3 26 105
use AOI22X1  AOI22X1_10
timestamp 1681708930
transform -1 0 1600 0 1 1970
box -8 -3 46 105
use NOR2X1  NOR2X1_21
timestamp 1681708930
transform -1 0 1624 0 1 1970
box -8 -3 32 105
use INVX2  INVX2_67
timestamp 1681708930
transform 1 0 1624 0 1 1970
box -9 -3 26 105
use M3_M2  M3_M2_828
timestamp 1681708930
transform 1 0 1692 0 1 1975
box -3 -3 3 3
use XNOR2X1  XNOR2X1_11
timestamp 1681708930
transform 1 0 1640 0 1 1970
box -8 -3 64 105
use FILL  FILL_341
timestamp 1681708930
transform 1 0 1696 0 1 1970
box -8 -3 16 105
use FILL  FILL_342
timestamp 1681708930
transform 1 0 1704 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_829
timestamp 1681708930
transform 1 0 1740 0 1 1975
box -3 -3 3 3
use NOR2X1  NOR2X1_22
timestamp 1681708930
transform 1 0 1712 0 1 1970
box -8 -3 32 105
use FILL  FILL_343
timestamp 1681708930
transform 1 0 1736 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_68
timestamp 1681708930
transform 1 0 1744 0 1 1970
box -9 -3 26 105
use FILL  FILL_344
timestamp 1681708930
transform 1 0 1760 0 1 1970
box -8 -3 16 105
use FILL  FILL_365
timestamp 1681708930
transform 1 0 1768 0 1 1970
box -8 -3 16 105
use NAND2X1  NAND2X1_35
timestamp 1681708930
transform -1 0 1800 0 1 1970
box -8 -3 32 105
use M3_M2  M3_M2_830
timestamp 1681708930
transform 1 0 1844 0 1 1975
box -3 -3 3 3
use AOI22X1  AOI22X1_11
timestamp 1681708930
transform 1 0 1800 0 1 1970
box -8 -3 46 105
use FILL  FILL_366
timestamp 1681708930
transform 1 0 1840 0 1 1970
box -8 -3 16 105
use FILL  FILL_367
timestamp 1681708930
transform 1 0 1848 0 1 1970
box -8 -3 16 105
use FILL  FILL_368
timestamp 1681708930
transform 1 0 1856 0 1 1970
box -8 -3 16 105
use FILL  FILL_369
timestamp 1681708930
transform 1 0 1864 0 1 1970
box -8 -3 16 105
use FILL  FILL_370
timestamp 1681708930
transform 1 0 1872 0 1 1970
box -8 -3 16 105
use FILL  FILL_371
timestamp 1681708930
transform 1 0 1880 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_831
timestamp 1681708930
transform 1 0 1908 0 1 1975
box -3 -3 3 3
use AOI22X1  AOI22X1_12
timestamp 1681708930
transform 1 0 1888 0 1 1970
box -8 -3 46 105
use FILL  FILL_372
timestamp 1681708930
transform 1 0 1928 0 1 1970
box -8 -3 16 105
use FILL  FILL_373
timestamp 1681708930
transform 1 0 1936 0 1 1970
box -8 -3 16 105
use FILL  FILL_374
timestamp 1681708930
transform 1 0 1944 0 1 1970
box -8 -3 16 105
use FILL  FILL_375
timestamp 1681708930
transform 1 0 1952 0 1 1970
box -8 -3 16 105
use FILL  FILL_376
timestamp 1681708930
transform 1 0 1960 0 1 1970
box -8 -3 16 105
use FILL  FILL_377
timestamp 1681708930
transform 1 0 1968 0 1 1970
box -8 -3 16 105
use FILL  FILL_378
timestamp 1681708930
transform 1 0 1976 0 1 1970
box -8 -3 16 105
use XOR2X1  XOR2X1_47
timestamp 1681708930
transform -1 0 2040 0 1 1970
box -8 -3 64 105
use INVX2  INVX2_72
timestamp 1681708930
transform -1 0 2056 0 1 1970
box -9 -3 26 105
use NOR2X1  NOR2X1_26
timestamp 1681708930
transform 1 0 2056 0 1 1970
box -8 -3 32 105
use FILL  FILL_379
timestamp 1681708930
transform 1 0 2080 0 1 1970
box -8 -3 16 105
use FILL  FILL_392
timestamp 1681708930
transform 1 0 2088 0 1 1970
box -8 -3 16 105
use FILL  FILL_393
timestamp 1681708930
transform 1 0 2096 0 1 1970
box -8 -3 16 105
use FILL  FILL_394
timestamp 1681708930
transform 1 0 2104 0 1 1970
box -8 -3 16 105
use FILL  FILL_396
timestamp 1681708930
transform 1 0 2112 0 1 1970
box -8 -3 16 105
use AOI21X1  AOI21X1_16
timestamp 1681708930
transform 1 0 2120 0 1 1970
box -7 -3 39 105
use FILL  FILL_397
timestamp 1681708930
transform 1 0 2152 0 1 1970
box -8 -3 16 105
use FILL  FILL_398
timestamp 1681708930
transform 1 0 2160 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_832
timestamp 1681708930
transform 1 0 2220 0 1 1975
box -3 -3 3 3
use XNOR2X1  XNOR2X1_13
timestamp 1681708930
transform -1 0 2224 0 1 1970
box -8 -3 64 105
use OAI21X1  OAI21X1_36
timestamp 1681708930
transform 1 0 2224 0 1 1970
box -8 -3 34 105
use FILL  FILL_399
timestamp 1681708930
transform 1 0 2256 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_833
timestamp 1681708930
transform 1 0 2284 0 1 1975
box -3 -3 3 3
use NAND2X1  NAND2X1_36
timestamp 1681708930
transform -1 0 2288 0 1 1970
box -8 -3 32 105
use FILL  FILL_400
timestamp 1681708930
transform 1 0 2288 0 1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_27
timestamp 1681708930
transform -1 0 2320 0 1 1970
box -8 -3 32 105
use FILL  FILL_401
timestamp 1681708930
transform 1 0 2320 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_13
timestamp 1681708930
transform -1 0 2368 0 1 1970
box -8 -3 46 105
use INVX2  INVX2_75
timestamp 1681708930
transform 1 0 2368 0 1 1970
box -9 -3 26 105
use XNOR2X1  XNOR2X1_14
timestamp 1681708930
transform 1 0 2384 0 1 1970
box -8 -3 64 105
use NAND2X1  NAND2X1_37
timestamp 1681708930
transform -1 0 2464 0 1 1970
box -8 -3 32 105
use OAI21X1  OAI21X1_37
timestamp 1681708930
transform 1 0 2464 0 1 1970
box -8 -3 34 105
use XOR2X1  XOR2X1_50
timestamp 1681708930
transform 1 0 2496 0 1 1970
box -8 -3 64 105
use XOR2X1  XOR2X1_51
timestamp 1681708930
transform 1 0 2552 0 1 1970
box -8 -3 64 105
use XOR2X1  XOR2X1_52
timestamp 1681708930
transform 1 0 2608 0 1 1970
box -8 -3 64 105
use top_mod_new_VIA0  top_mod_new_VIA0_13
timestamp 1681708930
transform 1 0 2688 0 1 1970
box -10 -3 10 3
use M3_M2  M3_M2_852
timestamp 1681708930
transform 1 0 76 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_876
timestamp 1681708930
transform 1 0 188 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_877
timestamp 1681708930
transform 1 0 228 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1009
timestamp 1681708930
transform 1 0 76 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1010
timestamp 1681708930
transform 1 0 124 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_895
timestamp 1681708930
transform 1 0 132 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_896
timestamp 1681708930
transform 1 0 164 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1011
timestamp 1681708930
transform 1 0 212 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1012
timestamp 1681708930
transform 1 0 228 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1076
timestamp 1681708930
transform 1 0 92 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_913
timestamp 1681708930
transform 1 0 124 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_1077
timestamp 1681708930
transform 1 0 132 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_914
timestamp 1681708930
transform 1 0 172 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_1078
timestamp 1681708930
transform 1 0 188 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_915
timestamp 1681708930
transform 1 0 228 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_853
timestamp 1681708930
transform 1 0 244 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_897
timestamp 1681708930
transform 1 0 236 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1013
timestamp 1681708930
transform 1 0 244 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_997
timestamp 1681708930
transform 1 0 260 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1014
timestamp 1681708930
transform 1 0 268 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1015
timestamp 1681708930
transform 1 0 276 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1079
timestamp 1681708930
transform 1 0 236 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_916
timestamp 1681708930
transform 1 0 252 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_1080
timestamp 1681708930
transform 1 0 260 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_932
timestamp 1681708930
transform 1 0 236 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_982
timestamp 1681708930
transform 1 0 260 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_878
timestamp 1681708930
transform 1 0 316 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1016
timestamp 1681708930
transform 1 0 316 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1081
timestamp 1681708930
transform 1 0 276 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1082
timestamp 1681708930
transform 1 0 284 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1083
timestamp 1681708930
transform 1 0 300 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_917
timestamp 1681708930
transform 1 0 308 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_1084
timestamp 1681708930
transform 1 0 316 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1085
timestamp 1681708930
transform 1 0 324 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_933
timestamp 1681708930
transform 1 0 284 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_934
timestamp 1681708930
transform 1 0 300 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_963
timestamp 1681708930
transform 1 0 276 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_964
timestamp 1681708930
transform 1 0 308 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_983
timestamp 1681708930
transform 1 0 292 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_854
timestamp 1681708930
transform 1 0 348 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_879
timestamp 1681708930
transform 1 0 332 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1017
timestamp 1681708930
transform 1 0 332 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1018
timestamp 1681708930
transform 1 0 340 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1086
timestamp 1681708930
transform 1 0 332 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_935
timestamp 1681708930
transform 1 0 332 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_834
timestamp 1681708930
transform 1 0 380 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_835
timestamp 1681708930
transform 1 0 404 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_836
timestamp 1681708930
transform 1 0 460 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_855
timestamp 1681708930
transform 1 0 396 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_1019
timestamp 1681708930
transform 1 0 364 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1020
timestamp 1681708930
transform 1 0 380 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1021
timestamp 1681708930
transform 1 0 468 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_918
timestamp 1681708930
transform 1 0 364 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_919
timestamp 1681708930
transform 1 0 380 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_1087
timestamp 1681708930
transform 1 0 404 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1088
timestamp 1681708930
transform 1 0 460 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1089
timestamp 1681708930
transform 1 0 476 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1142
timestamp 1681708930
transform 1 0 364 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_936
timestamp 1681708930
transform 1 0 404 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_965
timestamp 1681708930
transform 1 0 372 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_991
timestamp 1681708930
transform 1 0 348 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_992
timestamp 1681708930
transform 1 0 364 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_920
timestamp 1681708930
transform 1 0 484 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_1090
timestamp 1681708930
transform 1 0 492 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_856
timestamp 1681708930
transform 1 0 516 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_998
timestamp 1681708930
transform 1 0 516 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1022
timestamp 1681708930
transform 1 0 508 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1143
timestamp 1681708930
transform 1 0 484 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_937
timestamp 1681708930
transform 1 0 500 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_898
timestamp 1681708930
transform 1 0 524 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_837
timestamp 1681708930
transform 1 0 588 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_857
timestamp 1681708930
transform 1 0 572 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_999
timestamp 1681708930
transform 1 0 548 0 1 1945
box -2 -2 2 2
use M3_M2  M3_M2_880
timestamp 1681708930
transform 1 0 556 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_858
timestamp 1681708930
transform 1 0 644 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_881
timestamp 1681708930
transform 1 0 596 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_882
timestamp 1681708930
transform 1 0 612 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_883
timestamp 1681708930
transform 1 0 636 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1023
timestamp 1681708930
transform 1 0 540 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_899
timestamp 1681708930
transform 1 0 548 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1024
timestamp 1681708930
transform 1 0 572 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_900
timestamp 1681708930
transform 1 0 580 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1025
timestamp 1681708930
transform 1 0 596 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_901
timestamp 1681708930
transform 1 0 604 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1026
timestamp 1681708930
transform 1 0 612 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1091
timestamp 1681708930
transform 1 0 548 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1092
timestamp 1681708930
transform 1 0 556 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1093
timestamp 1681708930
transform 1 0 572 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1094
timestamp 1681708930
transform 1 0 588 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_938
timestamp 1681708930
transform 1 0 556 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_921
timestamp 1681708930
transform 1 0 596 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_902
timestamp 1681708930
transform 1 0 636 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1095
timestamp 1681708930
transform 1 0 604 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1096
timestamp 1681708930
transform 1 0 612 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_922
timestamp 1681708930
transform 1 0 620 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_939
timestamp 1681708930
transform 1 0 588 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_940
timestamp 1681708930
transform 1 0 612 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_1144
timestamp 1681708930
transform 1 0 644 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_838
timestamp 1681708930
transform 1 0 668 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_1027
timestamp 1681708930
transform 1 0 660 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1028
timestamp 1681708930
transform 1 0 668 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_941
timestamp 1681708930
transform 1 0 660 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_903
timestamp 1681708930
transform 1 0 684 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_859
timestamp 1681708930
transform 1 0 700 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_1000
timestamp 1681708930
transform 1 0 700 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1029
timestamp 1681708930
transform 1 0 692 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1097
timestamp 1681708930
transform 1 0 684 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_839
timestamp 1681708930
transform 1 0 716 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_1030
timestamp 1681708930
transform 1 0 716 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1098
timestamp 1681708930
transform 1 0 708 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_840
timestamp 1681708930
transform 1 0 764 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_860
timestamp 1681708930
transform 1 0 764 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_1001
timestamp 1681708930
transform 1 0 772 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1031
timestamp 1681708930
transform 1 0 764 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_923
timestamp 1681708930
transform 1 0 740 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_1099
timestamp 1681708930
transform 1 0 788 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_942
timestamp 1681708930
transform 1 0 788 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_841
timestamp 1681708930
transform 1 0 812 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_1032
timestamp 1681708930
transform 1 0 804 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1033
timestamp 1681708930
transform 1 0 812 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_861
timestamp 1681708930
transform 1 0 844 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_884
timestamp 1681708930
transform 1 0 836 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1034
timestamp 1681708930
transform 1 0 836 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1035
timestamp 1681708930
transform 1 0 844 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1100
timestamp 1681708930
transform 1 0 820 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_862
timestamp 1681708930
transform 1 0 956 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_885
timestamp 1681708930
transform 1 0 900 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1036
timestamp 1681708930
transform 1 0 876 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_904
timestamp 1681708930
transform 1 0 908 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_905
timestamp 1681708930
transform 1 0 924 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_886
timestamp 1681708930
transform 1 0 964 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1101
timestamp 1681708930
transform 1 0 900 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1102
timestamp 1681708930
transform 1 0 956 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1145
timestamp 1681708930
transform 1 0 860 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_966
timestamp 1681708930
transform 1 0 860 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_1037
timestamp 1681708930
transform 1 0 980 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_967
timestamp 1681708930
transform 1 0 972 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_842
timestamp 1681708930
transform 1 0 1012 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_843
timestamp 1681708930
transform 1 0 1036 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_844
timestamp 1681708930
transform 1 0 1108 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_845
timestamp 1681708930
transform 1 0 1148 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_846
timestamp 1681708930
transform 1 0 1236 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_863
timestamp 1681708930
transform 1 0 1100 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_887
timestamp 1681708930
transform 1 0 1028 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_888
timestamp 1681708930
transform 1 0 1092 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1038
timestamp 1681708930
transform 1 0 1012 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1039
timestamp 1681708930
transform 1 0 1100 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1103
timestamp 1681708930
transform 1 0 996 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1104
timestamp 1681708930
transform 1 0 1060 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1105
timestamp 1681708930
transform 1 0 1092 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1146
timestamp 1681708930
transform 1 0 996 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_968
timestamp 1681708930
transform 1 0 996 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_969
timestamp 1681708930
transform 1 0 1012 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_864
timestamp 1681708930
transform 1 0 1188 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_847
timestamp 1681708930
transform 1 0 1268 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_865
timestamp 1681708930
transform 1 0 1260 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_866
timestamp 1681708930
transform 1 0 1300 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_1040
timestamp 1681708930
transform 1 0 1148 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1041
timestamp 1681708930
transform 1 0 1164 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1042
timestamp 1681708930
transform 1 0 1252 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1681708930
transform 1 0 1148 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1107
timestamp 1681708930
transform 1 0 1204 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1108
timestamp 1681708930
transform 1 0 1244 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_943
timestamp 1681708930
transform 1 0 1148 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_924
timestamp 1681708930
transform 1 0 1252 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_970
timestamp 1681708930
transform 1 0 1164 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_971
timestamp 1681708930
transform 1 0 1212 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_1043
timestamp 1681708930
transform 1 0 1300 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1044
timestamp 1681708930
transform 1 0 1308 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_867
timestamp 1681708930
transform 1 0 1364 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_1045
timestamp 1681708930
transform 1 0 1356 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1046
timestamp 1681708930
transform 1 0 1364 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1109
timestamp 1681708930
transform 1 0 1308 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1110
timestamp 1681708930
transform 1 0 1332 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1111
timestamp 1681708930
transform 1 0 1340 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_944
timestamp 1681708930
transform 1 0 1308 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_945
timestamp 1681708930
transform 1 0 1340 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_1002
timestamp 1681708930
transform 1 0 1396 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1112
timestamp 1681708930
transform 1 0 1388 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_946
timestamp 1681708930
transform 1 0 1396 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_868
timestamp 1681708930
transform 1 0 1412 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_1113
timestamp 1681708930
transform 1 0 1412 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1114
timestamp 1681708930
transform 1 0 1436 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1115
timestamp 1681708930
transform 1 0 1460 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1047
timestamp 1681708930
transform 1 0 1484 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1147
timestamp 1681708930
transform 1 0 1508 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_925
timestamp 1681708930
transform 1 0 1532 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_1048
timestamp 1681708930
transform 1 0 1556 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1049
timestamp 1681708930
transform 1 0 1572 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1050
timestamp 1681708930
transform 1 0 1588 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1051
timestamp 1681708930
transform 1 0 1604 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1116
timestamp 1681708930
transform 1 0 1540 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1681708930
transform 1 0 1532 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_926
timestamp 1681708930
transform 1 0 1556 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_1117
timestamp 1681708930
transform 1 0 1564 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1681708930
transform 1 0 1580 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1119
timestamp 1681708930
transform 1 0 1596 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1120
timestamp 1681708930
transform 1 0 1604 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_947
timestamp 1681708930
transform 1 0 1564 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_948
timestamp 1681708930
transform 1 0 1596 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_1149
timestamp 1681708930
transform 1 0 1612 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_848
timestamp 1681708930
transform 1 0 1644 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_1052
timestamp 1681708930
transform 1 0 1636 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1053
timestamp 1681708930
transform 1 0 1644 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1121
timestamp 1681708930
transform 1 0 1636 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_927
timestamp 1681708930
transform 1 0 1652 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_1122
timestamp 1681708930
transform 1 0 1660 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_928
timestamp 1681708930
transform 1 0 1668 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_949
timestamp 1681708930
transform 1 0 1636 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_1054
timestamp 1681708930
transform 1 0 1692 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_906
timestamp 1681708930
transform 1 0 1700 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1123
timestamp 1681708930
transform 1 0 1692 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1124
timestamp 1681708930
transform 1 0 1700 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1150
timestamp 1681708930
transform 1 0 1684 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_950
timestamp 1681708930
transform 1 0 1692 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_1003
timestamp 1681708930
transform 1 0 1724 0 1 1945
box -2 -2 2 2
use M3_M2  M3_M2_907
timestamp 1681708930
transform 1 0 1732 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1055
timestamp 1681708930
transform 1 0 1740 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1125
timestamp 1681708930
transform 1 0 1724 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_929
timestamp 1681708930
transform 1 0 1732 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_1151
timestamp 1681708930
transform 1 0 1732 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1165
timestamp 1681708930
transform 1 0 1748 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_1056
timestamp 1681708930
transform 1 0 1788 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1152
timestamp 1681708930
transform 1 0 1780 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_993
timestamp 1681708930
transform 1 0 1796 0 1 1885
box -3 -3 3 3
use M2_M1  M2_M1_1004
timestamp 1681708930
transform 1 0 1820 0 1 1945
box -2 -2 2 2
use M3_M2  M3_M2_908
timestamp 1681708930
transform 1 0 1820 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1057
timestamp 1681708930
transform 1 0 1828 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_930
timestamp 1681708930
transform 1 0 1812 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_889
timestamp 1681708930
transform 1 0 1860 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_972
timestamp 1681708930
transform 1 0 1844 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_869
timestamp 1681708930
transform 1 0 1884 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_849
timestamp 1681708930
transform 1 0 1932 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_870
timestamp 1681708930
transform 1 0 1916 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_871
timestamp 1681708930
transform 1 0 1940 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_1058
timestamp 1681708930
transform 1 0 1884 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1059
timestamp 1681708930
transform 1 0 1908 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1060
timestamp 1681708930
transform 1 0 1924 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1126
timestamp 1681708930
transform 1 0 1868 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1127
timestamp 1681708930
transform 1 0 1916 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_931
timestamp 1681708930
transform 1 0 1924 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_872
timestamp 1681708930
transform 1 0 1988 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_1061
timestamp 1681708930
transform 1 0 1980 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_890
timestamp 1681708930
transform 1 0 2052 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1062
timestamp 1681708930
transform 1 0 2028 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1128
timestamp 1681708930
transform 1 0 1948 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1129
timestamp 1681708930
transform 1 0 1972 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1130
timestamp 1681708930
transform 1 0 2004 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1153
timestamp 1681708930
transform 1 0 1876 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_951
timestamp 1681708930
transform 1 0 1884 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_1154
timestamp 1681708930
transform 1 0 1900 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_952
timestamp 1681708930
transform 1 0 1908 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_1166
timestamp 1681708930
transform 1 0 1884 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_973
timestamp 1681708930
transform 1 0 1908 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_984
timestamp 1681708930
transform 1 0 1892 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_994
timestamp 1681708930
transform 1 0 1876 0 1 1885
box -3 -3 3 3
use M2_M1  M2_M1_1131
timestamp 1681708930
transform 1 0 2044 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1155
timestamp 1681708930
transform 1 0 2036 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_974
timestamp 1681708930
transform 1 0 2004 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_975
timestamp 1681708930
transform 1 0 2036 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_1167
timestamp 1681708930
transform 1 0 2052 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_985
timestamp 1681708930
transform 1 0 1972 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_986
timestamp 1681708930
transform 1 0 2020 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_987
timestamp 1681708930
transform 1 0 2044 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_995
timestamp 1681708930
transform 1 0 2012 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_996
timestamp 1681708930
transform 1 0 2028 0 1 1885
box -3 -3 3 3
use M2_M1  M2_M1_1063
timestamp 1681708930
transform 1 0 2076 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_953
timestamp 1681708930
transform 1 0 2076 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_988
timestamp 1681708930
transform 1 0 2068 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_997
timestamp 1681708930
transform 1 0 2076 0 1 1885
box -3 -3 3 3
use M2_M1  M2_M1_1156
timestamp 1681708930
transform 1 0 2084 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_909
timestamp 1681708930
transform 1 0 2100 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1132
timestamp 1681708930
transform 1 0 2100 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_850
timestamp 1681708930
transform 1 0 2132 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_873
timestamp 1681708930
transform 1 0 2156 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_1005
timestamp 1681708930
transform 1 0 2148 0 1 1945
box -2 -2 2 2
use M3_M2  M3_M2_910
timestamp 1681708930
transform 1 0 2148 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_851
timestamp 1681708930
transform 1 0 2172 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_891
timestamp 1681708930
transform 1 0 2164 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1064
timestamp 1681708930
transform 1 0 2156 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1065
timestamp 1681708930
transform 1 0 2164 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1133
timestamp 1681708930
transform 1 0 2124 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1157
timestamp 1681708930
transform 1 0 2116 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_954
timestamp 1681708930
transform 1 0 2124 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_1158
timestamp 1681708930
transform 1 0 2140 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1168
timestamp 1681708930
transform 1 0 2108 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_976
timestamp 1681708930
transform 1 0 2116 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_977
timestamp 1681708930
transform 1 0 2140 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_955
timestamp 1681708930
transform 1 0 2164 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_989
timestamp 1681708930
transform 1 0 2180 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_874
timestamp 1681708930
transform 1 0 2212 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_875
timestamp 1681708930
transform 1 0 2228 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_911
timestamp 1681708930
transform 1 0 2220 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1066
timestamp 1681708930
transform 1 0 2228 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1134
timestamp 1681708930
transform 1 0 2228 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1135
timestamp 1681708930
transform 1 0 2236 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1159
timestamp 1681708930
transform 1 0 2220 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_956
timestamp 1681708930
transform 1 0 2228 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_1160
timestamp 1681708930
transform 1 0 2244 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1161
timestamp 1681708930
transform 1 0 2252 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1067
timestamp 1681708930
transform 1 0 2260 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_978
timestamp 1681708930
transform 1 0 2252 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_990
timestamp 1681708930
transform 1 0 2244 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_1136
timestamp 1681708930
transform 1 0 2276 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_957
timestamp 1681708930
transform 1 0 2276 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_1068
timestamp 1681708930
transform 1 0 2292 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1069
timestamp 1681708930
transform 1 0 2316 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1137
timestamp 1681708930
transform 1 0 2324 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_892
timestamp 1681708930
transform 1 0 2348 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1070
timestamp 1681708930
transform 1 0 2348 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_893
timestamp 1681708930
transform 1 0 2388 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_912
timestamp 1681708930
transform 1 0 2388 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1071
timestamp 1681708930
transform 1 0 2396 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1072
timestamp 1681708930
transform 1 0 2404 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1138
timestamp 1681708930
transform 1 0 2380 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1139
timestamp 1681708930
transform 1 0 2396 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1162
timestamp 1681708930
transform 1 0 2364 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_958
timestamp 1681708930
transform 1 0 2388 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_1163
timestamp 1681708930
transform 1 0 2404 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_959
timestamp 1681708930
transform 1 0 2412 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_1006
timestamp 1681708930
transform 1 0 2428 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1007
timestamp 1681708930
transform 1 0 2436 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1164
timestamp 1681708930
transform 1 0 2420 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_979
timestamp 1681708930
transform 1 0 2404 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_1073
timestamp 1681708930
transform 1 0 2452 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1008
timestamp 1681708930
transform 1 0 2468 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1140
timestamp 1681708930
transform 1 0 2468 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_960
timestamp 1681708930
transform 1 0 2468 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_980
timestamp 1681708930
transform 1 0 2460 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_981
timestamp 1681708930
transform 1 0 2484 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_894
timestamp 1681708930
transform 1 0 2508 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1141
timestamp 1681708930
transform 1 0 2508 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_961
timestamp 1681708930
transform 1 0 2524 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_1074
timestamp 1681708930
transform 1 0 2532 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1075
timestamp 1681708930
transform 1 0 2540 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_962
timestamp 1681708930
transform 1 0 2596 0 1 1915
box -3 -3 3 3
use top_mod_new_VIA0  top_mod_new_VIA0_14
timestamp 1681708930
transform 1 0 24 0 1 1870
box -10 -3 10 3
use XNOR2X1  XNOR2X1_10
timestamp 1681708930
transform -1 0 128 0 -1 1970
box -8 -3 64 105
use DFFNEGX1  DFFNEGX1_26
timestamp 1681708930
transform -1 0 224 0 -1 1970
box -8 -3 104 105
use INVX2  INVX2_62
timestamp 1681708930
transform 1 0 224 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_63
timestamp 1681708930
transform 1 0 240 0 -1 1970
box -9 -3 26 105
use NOR2X1  NOR2X1_19
timestamp 1681708930
transform 1 0 256 0 -1 1970
box -8 -3 32 105
use AOI22X1  AOI22X1_8
timestamp 1681708930
transform 1 0 280 0 -1 1970
box -8 -3 46 105
use INVX2  INVX2_64
timestamp 1681708930
transform -1 0 336 0 -1 1970
box -9 -3 26 105
use OAI21X1  OAI21X1_31
timestamp 1681708930
transform 1 0 336 0 -1 1970
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_27
timestamp 1681708930
transform 1 0 368 0 -1 1970
box -8 -3 104 105
use NAND2X1  NAND2X1_27
timestamp 1681708930
transform 1 0 464 0 -1 1970
box -8 -3 32 105
use BUFX2  BUFX2_0
timestamp 1681708930
transform 1 0 488 0 -1 1970
box -5 -3 28 105
use FILL  FILL_332
timestamp 1681708930
transform 1 0 512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_333
timestamp 1681708930
transform 1 0 520 0 -1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_20
timestamp 1681708930
transform 1 0 528 0 -1 1970
box -8 -3 32 105
use M3_M2  M3_M2_998
timestamp 1681708930
transform 1 0 564 0 1 1875
box -3 -3 3 3
use INVX2  INVX2_65
timestamp 1681708930
transform 1 0 552 0 -1 1970
box -9 -3 26 105
use AOI22X1  AOI22X1_9
timestamp 1681708930
transform 1 0 568 0 -1 1970
box -8 -3 46 105
use OAI21X1  OAI21X1_32
timestamp 1681708930
transform 1 0 608 0 -1 1970
box -8 -3 34 105
use FILL  FILL_334
timestamp 1681708930
transform 1 0 640 0 -1 1970
box -8 -3 16 105
use FILL  FILL_336
timestamp 1681708930
transform 1 0 648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_345
timestamp 1681708930
transform 1 0 656 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_69
timestamp 1681708930
transform 1 0 664 0 -1 1970
box -9 -3 26 105
use NOR2X1  NOR2X1_23
timestamp 1681708930
transform -1 0 704 0 -1 1970
box -8 -3 32 105
use FILL  FILL_346
timestamp 1681708930
transform 1 0 704 0 -1 1970
box -8 -3 16 105
use XOR2X1  XOR2X1_44
timestamp 1681708930
transform -1 0 768 0 -1 1970
box -8 -3 64 105
use NOR2X1  NOR2X1_24
timestamp 1681708930
transform 1 0 768 0 -1 1970
box -8 -3 32 105
use FILL  FILL_347
timestamp 1681708930
transform 1 0 792 0 -1 1970
box -8 -3 16 105
use FILL  FILL_348
timestamp 1681708930
transform 1 0 800 0 -1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_34
timestamp 1681708930
transform 1 0 808 0 -1 1970
box -8 -3 34 105
use NAND2X1  NAND2X1_30
timestamp 1681708930
transform 1 0 840 0 -1 1970
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_31
timestamp 1681708930
transform 1 0 864 0 -1 1970
box -8 -3 104 105
use FILL  FILL_349
timestamp 1681708930
transform 1 0 960 0 -1 1970
box -8 -3 16 105
use FILL  FILL_350
timestamp 1681708930
transform 1 0 968 0 -1 1970
box -8 -3 16 105
use NAND2X1  NAND2X1_31
timestamp 1681708930
transform 1 0 976 0 -1 1970
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_32
timestamp 1681708930
transform 1 0 1000 0 -1 1970
box -8 -3 104 105
use XOR2X1  XOR2X1_45
timestamp 1681708930
transform 1 0 1096 0 -1 1970
box -8 -3 64 105
use DFFNEGX1  DFFNEGX1_33
timestamp 1681708930
transform 1 0 1152 0 -1 1970
box -8 -3 104 105
use M3_M2  M3_M2_999
timestamp 1681708930
transform 1 0 1308 0 1 1875
box -3 -3 3 3
use XNOR2X1  XNOR2X1_12
timestamp 1681708930
transform 1 0 1248 0 -1 1970
box -8 -3 64 105
use XOR2X1  XOR2X1_46
timestamp 1681708930
transform 1 0 1304 0 -1 1970
box -8 -3 64 105
use AOI21X1  AOI21X1_14
timestamp 1681708930
transform 1 0 1360 0 -1 1970
box -7 -3 39 105
use NOR2X1  NOR2X1_25
timestamp 1681708930
transform 1 0 1392 0 -1 1970
box -8 -3 32 105
use FILL  FILL_351
timestamp 1681708930
transform 1 0 1416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_352
timestamp 1681708930
transform 1 0 1424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_353
timestamp 1681708930
transform 1 0 1432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_354
timestamp 1681708930
transform 1 0 1440 0 -1 1970
box -8 -3 16 105
use FILL  FILL_355
timestamp 1681708930
transform 1 0 1448 0 -1 1970
box -8 -3 16 105
use FILL  FILL_356
timestamp 1681708930
transform 1 0 1456 0 -1 1970
box -8 -3 16 105
use FILL  FILL_357
timestamp 1681708930
transform 1 0 1464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_358
timestamp 1681708930
transform 1 0 1472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_359
timestamp 1681708930
transform 1 0 1480 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_1000
timestamp 1681708930
transform 1 0 1500 0 1 1875
box -3 -3 3 3
use NAND2X1  NAND2X1_32
timestamp 1681708930
transform 1 0 1488 0 -1 1970
box -8 -3 32 105
use FILL  FILL_360
timestamp 1681708930
transform 1 0 1512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_361
timestamp 1681708930
transform 1 0 1520 0 -1 1970
box -8 -3 16 105
use NAND2X1  NAND2X1_33
timestamp 1681708930
transform -1 0 1552 0 -1 1970
box -8 -3 32 105
use OAI22X1  OAI22X1_17
timestamp 1681708930
transform 1 0 1552 0 -1 1970
box -8 -3 46 105
use INVX2  INVX2_70
timestamp 1681708930
transform -1 0 1608 0 -1 1970
box -9 -3 26 105
use OAI21X1  OAI21X1_35
timestamp 1681708930
transform -1 0 1640 0 -1 1970
box -8 -3 34 105
use INVX2  INVX2_71
timestamp 1681708930
transform 1 0 1640 0 -1 1970
box -9 -3 26 105
use FILL  FILL_362
timestamp 1681708930
transform 1 0 1656 0 -1 1970
box -8 -3 16 105
use NAND2X1  NAND2X1_34
timestamp 1681708930
transform 1 0 1664 0 -1 1970
box -8 -3 32 105
use FILL  FILL_363
timestamp 1681708930
transform 1 0 1688 0 -1 1970
box -8 -3 16 105
use AOI21X1  AOI21X1_15
timestamp 1681708930
transform 1 0 1696 0 -1 1970
box -7 -3 39 105
use NAND3X1  NAND3X1_33
timestamp 1681708930
transform 1 0 1728 0 -1 1970
box -8 -3 40 105
use FILL  FILL_364
timestamp 1681708930
transform 1 0 1760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_380
timestamp 1681708930
transform 1 0 1768 0 -1 1970
box -8 -3 16 105
use FILL  FILL_381
timestamp 1681708930
transform 1 0 1776 0 -1 1970
box -8 -3 16 105
use FILL  FILL_382
timestamp 1681708930
transform 1 0 1784 0 -1 1970
box -8 -3 16 105
use FILL  FILL_383
timestamp 1681708930
transform 1 0 1792 0 -1 1970
box -8 -3 16 105
use FILL  FILL_384
timestamp 1681708930
transform 1 0 1800 0 -1 1970
box -8 -3 16 105
use FILL  FILL_385
timestamp 1681708930
transform 1 0 1808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_386
timestamp 1681708930
transform 1 0 1816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_387
timestamp 1681708930
transform 1 0 1824 0 -1 1970
box -8 -3 16 105
use FILL  FILL_388
timestamp 1681708930
transform 1 0 1832 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_1001
timestamp 1681708930
transform 1 0 1852 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1002
timestamp 1681708930
transform 1 0 1876 0 1 1875
box -3 -3 3 3
use OR2X1  OR2X1_6
timestamp 1681708930
transform 1 0 1840 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_34
timestamp 1681708930
transform 1 0 1872 0 -1 1970
box -8 -3 40 105
use INVX2  INVX2_73
timestamp 1681708930
transform 1 0 1904 0 -1 1970
box -9 -3 26 105
use XOR2X1  XOR2X1_48
timestamp 1681708930
transform 1 0 1920 0 -1 1970
box -8 -3 64 105
use XOR2X1  XOR2X1_49
timestamp 1681708930
transform -1 0 2032 0 -1 1970
box -8 -3 64 105
use NAND3X1  NAND3X1_35
timestamp 1681708930
transform 1 0 2032 0 -1 1970
box -8 -3 40 105
use FILL  FILL_389
timestamp 1681708930
transform 1 0 2064 0 -1 1970
box -8 -3 16 105
use FILL  FILL_390
timestamp 1681708930
transform 1 0 2072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_391
timestamp 1681708930
transform 1 0 2080 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_74
timestamp 1681708930
transform 1 0 2088 0 -1 1970
box -9 -3 26 105
use FILL  FILL_395
timestamp 1681708930
transform 1 0 2104 0 -1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_36
timestamp 1681708930
transform 1 0 2112 0 -1 1970
box -8 -3 40 105
use NOR2X1  NOR2X1_28
timestamp 1681708930
transform 1 0 2144 0 -1 1970
box -8 -3 32 105
use FILL  FILL_402
timestamp 1681708930
transform 1 0 2168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_403
timestamp 1681708930
transform 1 0 2176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_404
timestamp 1681708930
transform 1 0 2184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_405
timestamp 1681708930
transform 1 0 2192 0 -1 1970
box -8 -3 16 105
use NAND2X1  NAND2X1_38
timestamp 1681708930
transform 1 0 2200 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_39
timestamp 1681708930
transform 1 0 2224 0 -1 1970
box -8 -3 32 105
use FILL  FILL_406
timestamp 1681708930
transform 1 0 2248 0 -1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_38
timestamp 1681708930
transform -1 0 2288 0 -1 1970
box -8 -3 34 105
use FILL  FILL_407
timestamp 1681708930
transform 1 0 2288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_408
timestamp 1681708930
transform 1 0 2296 0 -1 1970
box -8 -3 16 105
use FILL  FILL_409
timestamp 1681708930
transform 1 0 2304 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_76
timestamp 1681708930
transform 1 0 2312 0 -1 1970
box -9 -3 26 105
use FILL  FILL_410
timestamp 1681708930
transform 1 0 2328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_411
timestamp 1681708930
transform 1 0 2336 0 -1 1970
box -8 -3 16 105
use NAND2X1  NAND2X1_40
timestamp 1681708930
transform 1 0 2344 0 -1 1970
box -8 -3 32 105
use OAI21X1  OAI21X1_39
timestamp 1681708930
transform 1 0 2368 0 -1 1970
box -8 -3 34 105
use NAND2X1  NAND2X1_41
timestamp 1681708930
transform 1 0 2400 0 -1 1970
box -8 -3 32 105
use FILL  FILL_412
timestamp 1681708930
transform 1 0 2424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_413
timestamp 1681708930
transform 1 0 2432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_414
timestamp 1681708930
transform 1 0 2440 0 -1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_29
timestamp 1681708930
transform 1 0 2448 0 -1 1970
box -8 -3 32 105
use FILL  FILL_415
timestamp 1681708930
transform 1 0 2472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_416
timestamp 1681708930
transform 1 0 2480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_417
timestamp 1681708930
transform 1 0 2488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_418
timestamp 1681708930
transform 1 0 2496 0 -1 1970
box -8 -3 16 105
use FILL  FILL_419
timestamp 1681708930
transform 1 0 2504 0 -1 1970
box -8 -3 16 105
use FILL  FILL_420
timestamp 1681708930
transform 1 0 2512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_421
timestamp 1681708930
transform 1 0 2520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_422
timestamp 1681708930
transform 1 0 2528 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_77
timestamp 1681708930
transform 1 0 2536 0 -1 1970
box -9 -3 26 105
use FILL  FILL_423
timestamp 1681708930
transform 1 0 2552 0 -1 1970
box -8 -3 16 105
use FILL  FILL_424
timestamp 1681708930
transform 1 0 2560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_425
timestamp 1681708930
transform 1 0 2568 0 -1 1970
box -8 -3 16 105
use FILL  FILL_426
timestamp 1681708930
transform 1 0 2576 0 -1 1970
box -8 -3 16 105
use FILL  FILL_427
timestamp 1681708930
transform 1 0 2584 0 -1 1970
box -8 -3 16 105
use FILL  FILL_428
timestamp 1681708930
transform 1 0 2592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_429
timestamp 1681708930
transform 1 0 2600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_430
timestamp 1681708930
transform 1 0 2608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_431
timestamp 1681708930
transform 1 0 2616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_432
timestamp 1681708930
transform 1 0 2624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_433
timestamp 1681708930
transform 1 0 2632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_434
timestamp 1681708930
transform 1 0 2640 0 -1 1970
box -8 -3 16 105
use FILL  FILL_435
timestamp 1681708930
transform 1 0 2648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_436
timestamp 1681708930
transform 1 0 2656 0 -1 1970
box -8 -3 16 105
use top_mod_new_VIA0  top_mod_new_VIA0_15
timestamp 1681708930
transform 1 0 2712 0 1 1870
box -10 -3 10 3
use M2_M1  M2_M1_1272
timestamp 1681708930
transform 1 0 92 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1025
timestamp 1681708930
transform 1 0 156 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1017
timestamp 1681708930
transform 1 0 180 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_1181
timestamp 1681708930
transform 1 0 156 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1210
timestamp 1681708930
transform 1 0 132 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1211
timestamp 1681708930
transform 1 0 148 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1043
timestamp 1681708930
transform 1 0 172 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_1273
timestamp 1681708930
transform 1 0 148 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1274
timestamp 1681708930
transform 1 0 156 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1275
timestamp 1681708930
transform 1 0 172 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1115
timestamp 1681708930
transform 1 0 140 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1116
timestamp 1681708930
transform 1 0 156 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_1182
timestamp 1681708930
transform 1 0 188 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1018
timestamp 1681708930
transform 1 0 220 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1026
timestamp 1681708930
transform 1 0 212 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_1183
timestamp 1681708930
transform 1 0 204 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1212
timestamp 1681708930
transform 1 0 196 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1276
timestamp 1681708930
transform 1 0 204 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1003
timestamp 1681708930
transform 1 0 244 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1019
timestamp 1681708930
transform 1 0 300 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1027
timestamp 1681708930
transform 1 0 284 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_1169
timestamp 1681708930
transform 1 0 292 0 1 1835
box -2 -2 2 2
use M3_M2  M3_M2_1028
timestamp 1681708930
transform 1 0 300 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_1184
timestamp 1681708930
transform 1 0 284 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1185
timestamp 1681708930
transform 1 0 300 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1073
timestamp 1681708930
transform 1 0 244 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1074
timestamp 1681708930
transform 1 0 260 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1213
timestamp 1681708930
transform 1 0 276 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1075
timestamp 1681708930
transform 1 0 284 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1277
timestamp 1681708930
transform 1 0 228 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1044
timestamp 1681708930
transform 1 0 316 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1076
timestamp 1681708930
transform 1 0 308 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1214
timestamp 1681708930
transform 1 0 316 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1278
timestamp 1681708930
transform 1 0 276 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1279
timestamp 1681708930
transform 1 0 300 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1132
timestamp 1681708930
transform 1 0 244 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1133
timestamp 1681708930
transform 1 0 260 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1117
timestamp 1681708930
transform 1 0 300 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1029
timestamp 1681708930
transform 1 0 332 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_1186
timestamp 1681708930
transform 1 0 348 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1077
timestamp 1681708930
transform 1 0 340 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1280
timestamp 1681708930
transform 1 0 340 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1004
timestamp 1681708930
transform 1 0 364 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1013
timestamp 1681708930
transform 1 0 372 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_1170
timestamp 1681708930
transform 1 0 364 0 1 1835
box -2 -2 2 2
use M3_M2  M3_M2_1030
timestamp 1681708930
transform 1 0 380 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_1187
timestamp 1681708930
transform 1 0 380 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1078
timestamp 1681708930
transform 1 0 364 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1215
timestamp 1681708930
transform 1 0 372 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1188
timestamp 1681708930
transform 1 0 396 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1216
timestamp 1681708930
transform 1 0 420 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1118
timestamp 1681708930
transform 1 0 404 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1134
timestamp 1681708930
transform 1 0 412 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1005
timestamp 1681708930
transform 1 0 452 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1006
timestamp 1681708930
transform 1 0 476 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1020
timestamp 1681708930
transform 1 0 460 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_1171
timestamp 1681708930
transform 1 0 452 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_1189
timestamp 1681708930
transform 1 0 444 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1281
timestamp 1681708930
transform 1 0 436 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1098
timestamp 1681708930
transform 1 0 444 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_1190
timestamp 1681708930
transform 1 0 468 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1217
timestamp 1681708930
transform 1 0 484 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1099
timestamp 1681708930
transform 1 0 492 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1119
timestamp 1681708930
transform 1 0 468 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1120
timestamp 1681708930
transform 1 0 500 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_1191
timestamp 1681708930
transform 1 0 508 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1021
timestamp 1681708930
transform 1 0 540 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_1172
timestamp 1681708930
transform 1 0 548 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_1192
timestamp 1681708930
transform 1 0 540 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1045
timestamp 1681708930
transform 1 0 548 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_1218
timestamp 1681708930
transform 1 0 540 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1282
timestamp 1681708930
transform 1 0 516 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1100
timestamp 1681708930
transform 1 0 524 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1135
timestamp 1681708930
transform 1 0 524 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_1219
timestamp 1681708930
transform 1 0 572 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1079
timestamp 1681708930
transform 1 0 580 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1283
timestamp 1681708930
transform 1 0 556 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1284
timestamp 1681708930
transform 1 0 604 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1285
timestamp 1681708930
transform 1 0 612 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1121
timestamp 1681708930
transform 1 0 604 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_1193
timestamp 1681708930
transform 1 0 636 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1080
timestamp 1681708930
transform 1 0 668 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1220
timestamp 1681708930
transform 1 0 676 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1221
timestamp 1681708930
transform 1 0 708 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1286
timestamp 1681708930
transform 1 0 636 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1287
timestamp 1681708930
transform 1 0 644 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1288
timestamp 1681708930
transform 1 0 652 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1289
timestamp 1681708930
transform 1 0 676 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1290
timestamp 1681708930
transform 1 0 684 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1136
timestamp 1681708930
transform 1 0 604 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1137
timestamp 1681708930
transform 1 0 628 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_1341
timestamp 1681708930
transform 1 0 668 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_1101
timestamp 1681708930
transform 1 0 700 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_1291
timestamp 1681708930
transform 1 0 708 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1342
timestamp 1681708930
transform 1 0 700 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_1138
timestamp 1681708930
transform 1 0 668 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1139
timestamp 1681708930
transform 1 0 692 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1140
timestamp 1681708930
transform 1 0 708 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1022
timestamp 1681708930
transform 1 0 732 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_1173
timestamp 1681708930
transform 1 0 724 0 1 1835
box -2 -2 2 2
use M3_M2  M3_M2_1046
timestamp 1681708930
transform 1 0 716 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_1194
timestamp 1681708930
transform 1 0 724 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1102
timestamp 1681708930
transform 1 0 748 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_1292
timestamp 1681708930
transform 1 0 756 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1195
timestamp 1681708930
transform 1 0 764 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1081
timestamp 1681708930
transform 1 0 764 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1047
timestamp 1681708930
transform 1 0 780 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_1222
timestamp 1681708930
transform 1 0 780 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1293
timestamp 1681708930
transform 1 0 772 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1082
timestamp 1681708930
transform 1 0 788 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1294
timestamp 1681708930
transform 1 0 788 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1083
timestamp 1681708930
transform 1 0 804 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1014
timestamp 1681708930
transform 1 0 820 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1084
timestamp 1681708930
transform 1 0 836 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1295
timestamp 1681708930
transform 1 0 836 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1223
timestamp 1681708930
transform 1 0 852 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1224
timestamp 1681708930
transform 1 0 916 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1296
timestamp 1681708930
transform 1 0 908 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1103
timestamp 1681708930
transform 1 0 916 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1007
timestamp 1681708930
transform 1 0 932 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1008
timestamp 1681708930
transform 1 0 1012 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1048
timestamp 1681708930
transform 1 0 980 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1049
timestamp 1681708930
transform 1 0 1020 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_1225
timestamp 1681708930
transform 1 0 980 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1226
timestamp 1681708930
transform 1 0 1012 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1227
timestamp 1681708930
transform 1 0 1020 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1297
timestamp 1681708930
transform 1 0 932 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1104
timestamp 1681708930
transform 1 0 996 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1105
timestamp 1681708930
transform 1 0 1012 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1141
timestamp 1681708930
transform 1 0 924 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_1298
timestamp 1681708930
transform 1 0 1044 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1228
timestamp 1681708930
transform 1 0 1060 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1106
timestamp 1681708930
transform 1 0 1060 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1142
timestamp 1681708930
transform 1 0 1084 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_1299
timestamp 1681708930
transform 1 0 1100 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1300
timestamp 1681708930
transform 1 0 1148 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1229
timestamp 1681708930
transform 1 0 1204 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1009
timestamp 1681708930
transform 1 0 1332 0 1 1865
box -3 -3 3 3
use M2_M1  M2_M1_1230
timestamp 1681708930
transform 1 0 1340 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1031
timestamp 1681708930
transform 1 0 1372 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_1196
timestamp 1681708930
transform 1 0 1372 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1174
timestamp 1681708930
transform 1 0 1412 0 1 1835
box -2 -2 2 2
use M3_M2  M3_M2_1010
timestamp 1681708930
transform 1 0 1484 0 1 1865
box -3 -3 3 3
use M2_M1  M2_M1_1197
timestamp 1681708930
transform 1 0 1412 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1231
timestamp 1681708930
transform 1 0 1404 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1050
timestamp 1681708930
transform 1 0 1444 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1051
timestamp 1681708930
transform 1 0 1476 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1052
timestamp 1681708930
transform 1 0 1492 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_1232
timestamp 1681708930
transform 1 0 1428 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1233
timestamp 1681708930
transform 1 0 1436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1234
timestamp 1681708930
transform 1 0 1452 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1085
timestamp 1681708930
transform 1 0 1460 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1235
timestamp 1681708930
transform 1 0 1468 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1236
timestamp 1681708930
transform 1 0 1476 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1237
timestamp 1681708930
transform 1 0 1492 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1238
timestamp 1681708930
transform 1 0 1508 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1301
timestamp 1681708930
transform 1 0 1420 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1302
timestamp 1681708930
transform 1 0 1436 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1303
timestamp 1681708930
transform 1 0 1444 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1304
timestamp 1681708930
transform 1 0 1460 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1122
timestamp 1681708930
transform 1 0 1420 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1123
timestamp 1681708930
transform 1 0 1436 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1143
timestamp 1681708930
transform 1 0 1428 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_1305
timestamp 1681708930
transform 1 0 1484 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1306
timestamp 1681708930
transform 1 0 1500 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1124
timestamp 1681708930
transform 1 0 1468 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1086
timestamp 1681708930
transform 1 0 1516 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1307
timestamp 1681708930
transform 1 0 1516 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1125
timestamp 1681708930
transform 1 0 1508 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_1343
timestamp 1681708930
transform 1 0 1516 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_1144
timestamp 1681708930
transform 1 0 1484 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1145
timestamp 1681708930
transform 1 0 1500 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1032
timestamp 1681708930
transform 1 0 1564 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_1175
timestamp 1681708930
transform 1 0 1572 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_1198
timestamp 1681708930
transform 1 0 1564 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1053
timestamp 1681708930
transform 1 0 1572 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_1239
timestamp 1681708930
transform 1 0 1556 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1240
timestamp 1681708930
transform 1 0 1572 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1199
timestamp 1681708930
transform 1 0 1596 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1054
timestamp 1681708930
transform 1 0 1644 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_1241
timestamp 1681708930
transform 1 0 1644 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1242
timestamp 1681708930
transform 1 0 1660 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1243
timestamp 1681708930
transform 1 0 1668 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1308
timestamp 1681708930
transform 1 0 1636 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1309
timestamp 1681708930
transform 1 0 1652 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1126
timestamp 1681708930
transform 1 0 1636 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1055
timestamp 1681708930
transform 1 0 1684 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_1310
timestamp 1681708930
transform 1 0 1676 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1311
timestamp 1681708930
transform 1 0 1684 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1056
timestamp 1681708930
transform 1 0 1732 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_1244
timestamp 1681708930
transform 1 0 1716 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1245
timestamp 1681708930
transform 1 0 1732 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1107
timestamp 1681708930
transform 1 0 1708 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_1344
timestamp 1681708930
transform 1 0 1708 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_1127
timestamp 1681708930
transform 1 0 1716 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_1312
timestamp 1681708930
transform 1 0 1748 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1128
timestamp 1681708930
transform 1 0 1748 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1087
timestamp 1681708930
transform 1 0 1780 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1246
timestamp 1681708930
transform 1 0 1796 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1313
timestamp 1681708930
transform 1 0 1780 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1314
timestamp 1681708930
transform 1 0 1788 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1108
timestamp 1681708930
transform 1 0 1796 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1129
timestamp 1681708930
transform 1 0 1788 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_1176
timestamp 1681708930
transform 1 0 1852 0 1 1835
box -2 -2 2 2
use M3_M2  M3_M2_1033
timestamp 1681708930
transform 1 0 1860 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_1200
timestamp 1681708930
transform 1 0 1836 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1201
timestamp 1681708930
transform 1 0 1844 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1247
timestamp 1681708930
transform 1 0 1820 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1057
timestamp 1681708930
transform 1 0 1852 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1058
timestamp 1681708930
transform 1 0 1868 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_1248
timestamp 1681708930
transform 1 0 1860 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1315
timestamp 1681708930
transform 1 0 1836 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1177
timestamp 1681708930
transform 1 0 1900 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_1178
timestamp 1681708930
transform 1 0 1908 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_1202
timestamp 1681708930
transform 1 0 1892 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1059
timestamp 1681708930
transform 1 0 1900 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1088
timestamp 1681708930
transform 1 0 1892 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1249
timestamp 1681708930
transform 1 0 1900 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1034
timestamp 1681708930
transform 1 0 1924 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_1203
timestamp 1681708930
transform 1 0 1932 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1060
timestamp 1681708930
transform 1 0 1940 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1061
timestamp 1681708930
transform 1 0 1980 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1089
timestamp 1681708930
transform 1 0 1972 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1316
timestamp 1681708930
transform 1 0 1948 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1090
timestamp 1681708930
transform 1 0 2004 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1317
timestamp 1681708930
transform 1 0 1996 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1023
timestamp 1681708930
transform 1 0 2020 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1035
timestamp 1681708930
transform 1 0 2052 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1062
timestamp 1681708930
transform 1 0 2036 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1063
timestamp 1681708930
transform 1 0 2060 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_1250
timestamp 1681708930
transform 1 0 2020 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1251
timestamp 1681708930
transform 1 0 2036 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1252
timestamp 1681708930
transform 1 0 2052 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1253
timestamp 1681708930
transform 1 0 2060 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1109
timestamp 1681708930
transform 1 0 2012 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_1318
timestamp 1681708930
transform 1 0 2028 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1146
timestamp 1681708930
transform 1 0 2020 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1011
timestamp 1681708930
transform 1 0 2092 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1091
timestamp 1681708930
transform 1 0 2076 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1015
timestamp 1681708930
transform 1 0 2108 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1024
timestamp 1681708930
transform 1 0 2108 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_1179
timestamp 1681708930
transform 1 0 2116 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_1204
timestamp 1681708930
transform 1 0 2100 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1205
timestamp 1681708930
transform 1 0 2108 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1206
timestamp 1681708930
transform 1 0 2132 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1319
timestamp 1681708930
transform 1 0 2068 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1320
timestamp 1681708930
transform 1 0 2076 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1147
timestamp 1681708930
transform 1 0 2060 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1110
timestamp 1681708930
transform 1 0 2084 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1092
timestamp 1681708930
transform 1 0 2116 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1321
timestamp 1681708930
transform 1 0 2100 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1322
timestamp 1681708930
transform 1 0 2116 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1323
timestamp 1681708930
transform 1 0 2140 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1130
timestamp 1681708930
transform 1 0 2100 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1148
timestamp 1681708930
transform 1 0 2092 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_1345
timestamp 1681708930
transform 1 0 2140 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_1149
timestamp 1681708930
transform 1 0 2140 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1036
timestamp 1681708930
transform 1 0 2188 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1064
timestamp 1681708930
transform 1 0 2172 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_1207
timestamp 1681708930
transform 1 0 2188 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1012
timestamp 1681708930
transform 1 0 2204 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1016
timestamp 1681708930
transform 1 0 2212 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_1254
timestamp 1681708930
transform 1 0 2164 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1255
timestamp 1681708930
transform 1 0 2172 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1256
timestamp 1681708930
transform 1 0 2188 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1093
timestamp 1681708930
transform 1 0 2196 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1324
timestamp 1681708930
transform 1 0 2156 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1111
timestamp 1681708930
transform 1 0 2172 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1065
timestamp 1681708930
transform 1 0 2228 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1066
timestamp 1681708930
transform 1 0 2260 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_1257
timestamp 1681708930
transform 1 0 2228 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1258
timestamp 1681708930
transform 1 0 2260 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1325
timestamp 1681708930
transform 1 0 2188 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1326
timestamp 1681708930
transform 1 0 2196 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1327
timestamp 1681708930
transform 1 0 2212 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1150
timestamp 1681708930
transform 1 0 2180 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_1259
timestamp 1681708930
transform 1 0 2292 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1328
timestamp 1681708930
transform 1 0 2260 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1329
timestamp 1681708930
transform 1 0 2276 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1151
timestamp 1681708930
transform 1 0 2260 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_1330
timestamp 1681708930
transform 1 0 2300 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1346
timestamp 1681708930
transform 1 0 2292 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_1131
timestamp 1681708930
transform 1 0 2300 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1067
timestamp 1681708930
transform 1 0 2340 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_1260
timestamp 1681708930
transform 1 0 2332 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1261
timestamp 1681708930
transform 1 0 2340 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1037
timestamp 1681708930
transform 1 0 2372 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1038
timestamp 1681708930
transform 1 0 2420 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1068
timestamp 1681708930
transform 1 0 2404 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1094
timestamp 1681708930
transform 1 0 2388 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1262
timestamp 1681708930
transform 1 0 2404 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1263
timestamp 1681708930
transform 1 0 2420 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1331
timestamp 1681708930
transform 1 0 2348 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1332
timestamp 1681708930
transform 1 0 2364 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1333
timestamp 1681708930
transform 1 0 2372 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1347
timestamp 1681708930
transform 1 0 2364 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_1095
timestamp 1681708930
transform 1 0 2428 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1334
timestamp 1681708930
transform 1 0 2428 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1152
timestamp 1681708930
transform 1 0 2428 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_1264
timestamp 1681708930
transform 1 0 2444 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1265
timestamp 1681708930
transform 1 0 2452 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1335
timestamp 1681708930
transform 1 0 2460 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1112
timestamp 1681708930
transform 1 0 2468 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_1208
timestamp 1681708930
transform 1 0 2484 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1266
timestamp 1681708930
transform 1 0 2484 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1348
timestamp 1681708930
transform 1 0 2476 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_1039
timestamp 1681708930
transform 1 0 2492 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1153
timestamp 1681708930
transform 1 0 2500 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_1180
timestamp 1681708930
transform 1 0 2532 0 1 1835
box -2 -2 2 2
use M3_M2  M3_M2_1040
timestamp 1681708930
transform 1 0 2548 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1069
timestamp 1681708930
transform 1 0 2540 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_1209
timestamp 1681708930
transform 1 0 2548 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1096
timestamp 1681708930
transform 1 0 2532 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1267
timestamp 1681708930
transform 1 0 2540 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1113
timestamp 1681708930
transform 1 0 2548 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1041
timestamp 1681708930
transform 1 0 2596 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1042
timestamp 1681708930
transform 1 0 2620 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1070
timestamp 1681708930
transform 1 0 2588 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1071
timestamp 1681708930
transform 1 0 2604 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_1268
timestamp 1681708930
transform 1 0 2580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1269
timestamp 1681708930
transform 1 0 2596 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1097
timestamp 1681708930
transform 1 0 2604 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_1270
timestamp 1681708930
transform 1 0 2620 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1271
timestamp 1681708930
transform 1 0 2628 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1336
timestamp 1681708930
transform 1 0 2564 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1337
timestamp 1681708930
transform 1 0 2572 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1338
timestamp 1681708930
transform 1 0 2588 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1114
timestamp 1681708930
transform 1 0 2596 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_1339
timestamp 1681708930
transform 1 0 2604 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1349
timestamp 1681708930
transform 1 0 2604 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_1340
timestamp 1681708930
transform 1 0 2620 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1154
timestamp 1681708930
transform 1 0 2572 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1155
timestamp 1681708930
transform 1 0 2604 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1156
timestamp 1681708930
transform 1 0 2628 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1072
timestamp 1681708930
transform 1 0 2644 0 1 1825
box -3 -3 3 3
use top_mod_new_VIA0  top_mod_new_VIA0_16
timestamp 1681708930
transform 1 0 48 0 1 1770
box -10 -3 10 3
use FILL  FILL_437
timestamp 1681708930
transform 1 0 72 0 1 1770
box -8 -3 16 105
use FILL  FILL_439
timestamp 1681708930
transform 1 0 80 0 1 1770
box -8 -3 16 105
use FILL  FILL_441
timestamp 1681708930
transform 1 0 88 0 1 1770
box -8 -3 16 105
use FILL  FILL_442
timestamp 1681708930
transform 1 0 96 0 1 1770
box -8 -3 16 105
use FILL  FILL_443
timestamp 1681708930
transform 1 0 104 0 1 1770
box -8 -3 16 105
use FILL  FILL_444
timestamp 1681708930
transform 1 0 112 0 1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_40
timestamp 1681708930
transform 1 0 120 0 1 1770
box -8 -3 34 105
use NAND2X1  NAND2X1_42
timestamp 1681708930
transform 1 0 152 0 1 1770
box -8 -3 32 105
use FILL  FILL_446
timestamp 1681708930
transform 1 0 176 0 1 1770
box -8 -3 16 105
use NAND2X1  NAND2X1_43
timestamp 1681708930
transform 1 0 184 0 1 1770
box -8 -3 32 105
use FILL  FILL_447
timestamp 1681708930
transform 1 0 208 0 1 1770
box -8 -3 16 105
use FILL  FILL_448
timestamp 1681708930
transform 1 0 216 0 1 1770
box -8 -3 16 105
use XNOR2X1  XNOR2X1_15
timestamp 1681708930
transform 1 0 224 0 1 1770
box -8 -3 64 105
use NAND3X1  NAND3X1_37
timestamp 1681708930
transform -1 0 312 0 1 1770
box -8 -3 40 105
use NOR2X1  NOR2X1_31
timestamp 1681708930
transform -1 0 336 0 1 1770
box -8 -3 32 105
use FILL  FILL_449
timestamp 1681708930
transform 1 0 336 0 1 1770
box -8 -3 16 105
use FILL  FILL_458
timestamp 1681708930
transform 1 0 344 0 1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_38
timestamp 1681708930
transform -1 0 384 0 1 1770
box -8 -3 40 105
use FILL  FILL_459
timestamp 1681708930
transform 1 0 384 0 1 1770
box -8 -3 16 105
use FILL  FILL_463
timestamp 1681708930
transform 1 0 392 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_1157
timestamp 1681708930
transform 1 0 436 0 1 1775
box -3 -3 3 3
use NAND3X1  NAND3X1_39
timestamp 1681708930
transform -1 0 432 0 1 1770
box -8 -3 40 105
use FILL  FILL_464
timestamp 1681708930
transform 1 0 432 0 1 1770
box -8 -3 16 105
use FILL  FILL_465
timestamp 1681708930
transform 1 0 440 0 1 1770
box -8 -3 16 105
use NAND2X1  NAND2X1_45
timestamp 1681708930
transform 1 0 448 0 1 1770
box -8 -3 32 105
use OAI21X1  OAI21X1_43
timestamp 1681708930
transform 1 0 472 0 1 1770
box -8 -3 34 105
use FILL  FILL_466
timestamp 1681708930
transform 1 0 504 0 1 1770
box -8 -3 16 105
use FILL  FILL_468
timestamp 1681708930
transform 1 0 512 0 1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_40
timestamp 1681708930
transform -1 0 552 0 1 1770
box -8 -3 40 105
use M3_M2  M3_M2_1158
timestamp 1681708930
transform 1 0 588 0 1 1775
box -3 -3 3 3
use XNOR2X1  XNOR2X1_17
timestamp 1681708930
transform -1 0 608 0 1 1770
box -8 -3 64 105
use OAI21X1  OAI21X1_45
timestamp 1681708930
transform 1 0 608 0 1 1770
box -8 -3 34 105
use AOI21X1  AOI21X1_18
timestamp 1681708930
transform 1 0 640 0 1 1770
box -7 -3 39 105
use M3_M2  M3_M2_1159
timestamp 1681708930
transform 1 0 684 0 1 1775
box -3 -3 3 3
use AOI21X1  AOI21X1_19
timestamp 1681708930
transform 1 0 672 0 1 1770
box -7 -3 39 105
use INVX2  INVX2_79
timestamp 1681708930
transform 1 0 704 0 1 1770
box -9 -3 26 105
use NAND3X1  NAND3X1_41
timestamp 1681708930
transform 1 0 720 0 1 1770
box -8 -3 40 105
use FILL  FILL_469
timestamp 1681708930
transform 1 0 752 0 1 1770
box -8 -3 16 105
use FILL  FILL_470
timestamp 1681708930
transform 1 0 760 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_80
timestamp 1681708930
transform 1 0 768 0 1 1770
box -9 -3 26 105
use FILL  FILL_471
timestamp 1681708930
transform 1 0 784 0 1 1770
box -8 -3 16 105
use FILL  FILL_483
timestamp 1681708930
transform 1 0 792 0 1 1770
box -8 -3 16 105
use FILL  FILL_485
timestamp 1681708930
transform 1 0 800 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_1160
timestamp 1681708930
transform 1 0 820 0 1 1775
box -3 -3 3 3
use FILL  FILL_486
timestamp 1681708930
transform 1 0 808 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_82
timestamp 1681708930
transform 1 0 816 0 1 1770
box -9 -3 26 105
use FILL  FILL_487
timestamp 1681708930
transform 1 0 832 0 1 1770
box -8 -3 16 105
use FILL  FILL_488
timestamp 1681708930
transform 1 0 840 0 1 1770
box -8 -3 16 105
use FILL  FILL_489
timestamp 1681708930
transform 1 0 848 0 1 1770
box -8 -3 16 105
use XNOR2X1  XNOR2X1_18
timestamp 1681708930
transform 1 0 856 0 1 1770
box -8 -3 64 105
use FILL  FILL_490
timestamp 1681708930
transform 1 0 912 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_1161
timestamp 1681708930
transform 1 0 948 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1162
timestamp 1681708930
transform 1 0 964 0 1 1775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_34
timestamp 1681708930
transform 1 0 920 0 1 1770
box -8 -3 104 105
use INVX2  INVX2_83
timestamp 1681708930
transform -1 0 1032 0 1 1770
box -9 -3 26 105
use FILL  FILL_492
timestamp 1681708930
transform 1 0 1032 0 1 1770
box -8 -3 16 105
use FILL  FILL_493
timestamp 1681708930
transform 1 0 1040 0 1 1770
box -8 -3 16 105
use FILL  FILL_494
timestamp 1681708930
transform 1 0 1048 0 1 1770
box -8 -3 16 105
use FILL  FILL_495
timestamp 1681708930
transform 1 0 1056 0 1 1770
box -8 -3 16 105
use FILL  FILL_496
timestamp 1681708930
transform 1 0 1064 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_84
timestamp 1681708930
transform -1 0 1088 0 1 1770
box -9 -3 26 105
use FILL  FILL_497
timestamp 1681708930
transform 1 0 1088 0 1 1770
box -8 -3 16 105
use FILL  FILL_498
timestamp 1681708930
transform 1 0 1096 0 1 1770
box -8 -3 16 105
use FILL  FILL_499
timestamp 1681708930
transform 1 0 1104 0 1 1770
box -8 -3 16 105
use FILL  FILL_500
timestamp 1681708930
transform 1 0 1112 0 1 1770
box -8 -3 16 105
use FILL  FILL_501
timestamp 1681708930
transform 1 0 1120 0 1 1770
box -8 -3 16 105
use FILL  FILL_511
timestamp 1681708930
transform 1 0 1128 0 1 1770
box -8 -3 16 105
use FILL  FILL_512
timestamp 1681708930
transform 1 0 1136 0 1 1770
box -8 -3 16 105
use FILL  FILL_513
timestamp 1681708930
transform 1 0 1144 0 1 1770
box -8 -3 16 105
use FILL  FILL_514
timestamp 1681708930
transform 1 0 1152 0 1 1770
box -8 -3 16 105
use FILL  FILL_515
timestamp 1681708930
transform 1 0 1160 0 1 1770
box -8 -3 16 105
use FILL  FILL_516
timestamp 1681708930
transform 1 0 1168 0 1 1770
box -8 -3 16 105
use FILL  FILL_517
timestamp 1681708930
transform 1 0 1176 0 1 1770
box -8 -3 16 105
use FILL  FILL_518
timestamp 1681708930
transform 1 0 1184 0 1 1770
box -8 -3 16 105
use FILL  FILL_520
timestamp 1681708930
transform 1 0 1192 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_86
timestamp 1681708930
transform 1 0 1200 0 1 1770
box -9 -3 26 105
use FILL  FILL_522
timestamp 1681708930
transform 1 0 1216 0 1 1770
box -8 -3 16 105
use FILL  FILL_523
timestamp 1681708930
transform 1 0 1224 0 1 1770
box -8 -3 16 105
use FILL  FILL_524
timestamp 1681708930
transform 1 0 1232 0 1 1770
box -8 -3 16 105
use FILL  FILL_525
timestamp 1681708930
transform 1 0 1240 0 1 1770
box -8 -3 16 105
use FILL  FILL_526
timestamp 1681708930
transform 1 0 1248 0 1 1770
box -8 -3 16 105
use FILL  FILL_527
timestamp 1681708930
transform 1 0 1256 0 1 1770
box -8 -3 16 105
use FILL  FILL_528
timestamp 1681708930
transform 1 0 1264 0 1 1770
box -8 -3 16 105
use FILL  FILL_529
timestamp 1681708930
transform 1 0 1272 0 1 1770
box -8 -3 16 105
use FILL  FILL_530
timestamp 1681708930
transform 1 0 1280 0 1 1770
box -8 -3 16 105
use FILL  FILL_531
timestamp 1681708930
transform 1 0 1288 0 1 1770
box -8 -3 16 105
use FILL  FILL_532
timestamp 1681708930
transform 1 0 1296 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_87
timestamp 1681708930
transform -1 0 1320 0 1 1770
box -9 -3 26 105
use FILL  FILL_533
timestamp 1681708930
transform 1 0 1320 0 1 1770
box -8 -3 16 105
use FILL  FILL_534
timestamp 1681708930
transform 1 0 1328 0 1 1770
box -8 -3 16 105
use FILL  FILL_535
timestamp 1681708930
transform 1 0 1336 0 1 1770
box -8 -3 16 105
use FILL  FILL_536
timestamp 1681708930
transform 1 0 1344 0 1 1770
box -8 -3 16 105
use FILL  FILL_537
timestamp 1681708930
transform 1 0 1352 0 1 1770
box -8 -3 16 105
use FILL  FILL_538
timestamp 1681708930
transform 1 0 1360 0 1 1770
box -8 -3 16 105
use FILL  FILL_539
timestamp 1681708930
transform 1 0 1368 0 1 1770
box -8 -3 16 105
use FILL  FILL_540
timestamp 1681708930
transform 1 0 1376 0 1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_45
timestamp 1681708930
transform -1 0 1416 0 1 1770
box -8 -3 40 105
use INVX2  INVX2_88
timestamp 1681708930
transform 1 0 1416 0 1 1770
box -9 -3 26 105
use AOI22X1  AOI22X1_18
timestamp 1681708930
transform 1 0 1432 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_19
timestamp 1681708930
transform 1 0 1472 0 1 1770
box -8 -3 46 105
use M3_M2  M3_M2_1163
timestamp 1681708930
transform 1 0 1524 0 1 1775
box -3 -3 3 3
use FILL  FILL_541
timestamp 1681708930
transform 1 0 1512 0 1 1770
box -8 -3 16 105
use FILL  FILL_542
timestamp 1681708930
transform 1 0 1520 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_1164
timestamp 1681708930
transform 1 0 1556 0 1 1775
box -3 -3 3 3
use OR2X1  OR2X1_7
timestamp 1681708930
transform 1 0 1528 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_46
timestamp 1681708930
transform 1 0 1560 0 1 1770
box -8 -3 40 105
use FILL  FILL_543
timestamp 1681708930
transform 1 0 1592 0 1 1770
box -8 -3 16 105
use FILL  FILL_544
timestamp 1681708930
transform 1 0 1600 0 1 1770
box -8 -3 16 105
use FILL  FILL_545
timestamp 1681708930
transform 1 0 1608 0 1 1770
box -8 -3 16 105
use FILL  FILL_546
timestamp 1681708930
transform 1 0 1616 0 1 1770
box -8 -3 16 105
use FILL  FILL_547
timestamp 1681708930
transform 1 0 1624 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_19
timestamp 1681708930
transform -1 0 1672 0 1 1770
box -8 -3 46 105
use FILL  FILL_548
timestamp 1681708930
transform 1 0 1672 0 1 1770
box -8 -3 16 105
use FILL  FILL_549
timestamp 1681708930
transform 1 0 1680 0 1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_37
timestamp 1681708930
transform -1 0 1712 0 1 1770
box -8 -3 32 105
use AOI22X1  AOI22X1_20
timestamp 1681708930
transform 1 0 1712 0 1 1770
box -8 -3 46 105
use FILL  FILL_550
timestamp 1681708930
transform 1 0 1752 0 1 1770
box -8 -3 16 105
use FILL  FILL_551
timestamp 1681708930
transform 1 0 1760 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_91
timestamp 1681708930
transform -1 0 1784 0 1 1770
box -9 -3 26 105
use FILL  FILL_552
timestamp 1681708930
transform 1 0 1784 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_92
timestamp 1681708930
transform 1 0 1792 0 1 1770
box -9 -3 26 105
use OAI21X1  OAI21X1_46
timestamp 1681708930
transform 1 0 1808 0 1 1770
box -8 -3 34 105
use NAND3X1  NAND3X1_47
timestamp 1681708930
transform -1 0 1872 0 1 1770
box -8 -3 40 105
use FILL  FILL_553
timestamp 1681708930
transform 1 0 1872 0 1 1770
box -8 -3 16 105
use FILL  FILL_554
timestamp 1681708930
transform 1 0 1880 0 1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_48
timestamp 1681708930
transform 1 0 1888 0 1 1770
box -8 -3 40 105
use FILL  FILL_555
timestamp 1681708930
transform 1 0 1920 0 1 1770
box -8 -3 16 105
use FILL  FILL_556
timestamp 1681708930
transform 1 0 1928 0 1 1770
box -8 -3 16 105
use FILL  FILL_565
timestamp 1681708930
transform 1 0 1936 0 1 1770
box -8 -3 16 105
use XOR2X1  XOR2X1_60
timestamp 1681708930
transform 1 0 1944 0 1 1770
box -8 -3 64 105
use FILL  FILL_566
timestamp 1681708930
transform 1 0 2000 0 1 1770
box -8 -3 16 105
use FILL  FILL_567
timestamp 1681708930
transform 1 0 2008 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_21
timestamp 1681708930
transform -1 0 2056 0 1 1770
box -8 -3 46 105
use FILL  FILL_568
timestamp 1681708930
transform 1 0 2056 0 1 1770
box -8 -3 16 105
use FILL  FILL_569
timestamp 1681708930
transform 1 0 2064 0 1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_48
timestamp 1681708930
transform 1 0 2072 0 1 1770
box -8 -3 34 105
use M3_M2  M3_M2_1165
timestamp 1681708930
transform 1 0 2116 0 1 1775
box -3 -3 3 3
use NAND3X1  NAND3X1_50
timestamp 1681708930
transform 1 0 2104 0 1 1770
box -8 -3 40 105
use M3_M2  M3_M2_1166
timestamp 1681708930
transform 1 0 2156 0 1 1775
box -3 -3 3 3
use NOR2X1  NOR2X1_38
timestamp 1681708930
transform 1 0 2136 0 1 1770
box -8 -3 32 105
use OAI21X1  OAI21X1_49
timestamp 1681708930
transform 1 0 2160 0 1 1770
box -8 -3 34 105
use INVX2  INVX2_95
timestamp 1681708930
transform 1 0 2192 0 1 1770
box -9 -3 26 105
use XNOR2X1  XNOR2X1_21
timestamp 1681708930
transform -1 0 2264 0 1 1770
box -8 -3 64 105
use AOI21X1  AOI21X1_22
timestamp 1681708930
transform 1 0 2264 0 1 1770
box -7 -3 39 105
use FILL  FILL_575
timestamp 1681708930
transform 1 0 2296 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_1167
timestamp 1681708930
transform 1 0 2348 0 1 1775
box -3 -3 3 3
use OR2X1  OR2X1_8
timestamp 1681708930
transform 1 0 2304 0 1 1770
box -8 -3 40 105
use M3_M2  M3_M2_1168
timestamp 1681708930
transform 1 0 2364 0 1 1775
box -3 -3 3 3
use AOI21X1  AOI21X1_23
timestamp 1681708930
transform 1 0 2336 0 1 1770
box -7 -3 39 105
use M3_M2  M3_M2_1169
timestamp 1681708930
transform 1 0 2388 0 1 1775
box -3 -3 3 3
use XNOR2X1  XNOR2X1_22
timestamp 1681708930
transform 1 0 2368 0 1 1770
box -8 -3 64 105
use M3_M2  M3_M2_1170
timestamp 1681708930
transform 1 0 2436 0 1 1775
box -3 -3 3 3
use FILL  FILL_576
timestamp 1681708930
transform 1 0 2424 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_96
timestamp 1681708930
transform -1 0 2448 0 1 1770
box -9 -3 26 105
use AOI21X1  AOI21X1_24
timestamp 1681708930
transform 1 0 2448 0 1 1770
box -7 -3 39 105
use FILL  FILL_577
timestamp 1681708930
transform 1 0 2480 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_1171
timestamp 1681708930
transform 1 0 2500 0 1 1775
box -3 -3 3 3
use FILL  FILL_578
timestamp 1681708930
transform 1 0 2488 0 1 1770
box -8 -3 16 105
use FILL  FILL_579
timestamp 1681708930
transform 1 0 2496 0 1 1770
box -8 -3 16 105
use FILL  FILL_580
timestamp 1681708930
transform 1 0 2504 0 1 1770
box -8 -3 16 105
use FILL  FILL_581
timestamp 1681708930
transform 1 0 2512 0 1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_51
timestamp 1681708930
transform -1 0 2552 0 1 1770
box -8 -3 40 105
use FILL  FILL_582
timestamp 1681708930
transform 1 0 2552 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_22
timestamp 1681708930
transform 1 0 2560 0 1 1770
box -8 -3 46 105
use M3_M2  M3_M2_1172
timestamp 1681708930
transform 1 0 2620 0 1 1775
box -3 -3 3 3
use NOR2X1  NOR2X1_39
timestamp 1681708930
transform 1 0 2600 0 1 1770
box -8 -3 32 105
use FILL  FILL_583
timestamp 1681708930
transform 1 0 2624 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_97
timestamp 1681708930
transform 1 0 2632 0 1 1770
box -9 -3 26 105
use FILL  FILL_584
timestamp 1681708930
transform 1 0 2648 0 1 1770
box -8 -3 16 105
use FILL  FILL_597
timestamp 1681708930
transform 1 0 2656 0 1 1770
box -8 -3 16 105
use top_mod_new_VIA0  top_mod_new_VIA0_17
timestamp 1681708930
transform 1 0 2688 0 1 1770
box -10 -3 10 3
use M2_M1  M2_M1_1350
timestamp 1681708930
transform 1 0 76 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1351
timestamp 1681708930
transform 1 0 92 0 1 1745
box -2 -2 2 2
use M3_M2  M3_M2_1200
timestamp 1681708930
transform 1 0 108 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_1363
timestamp 1681708930
transform 1 0 100 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1364
timestamp 1681708930
transform 1 0 108 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1437
timestamp 1681708930
transform 1 0 124 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1286
timestamp 1681708930
transform 1 0 124 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_1503
timestamp 1681708930
transform 1 0 140 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_1287
timestamp 1681708930
transform 1 0 140 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1201
timestamp 1681708930
transform 1 0 164 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1181
timestamp 1681708930
transform 1 0 196 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1182
timestamp 1681708930
transform 1 0 220 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_1352
timestamp 1681708930
transform 1 0 180 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1365
timestamp 1681708930
transform 1 0 164 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1366
timestamp 1681708930
transform 1 0 172 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1367
timestamp 1681708930
transform 1 0 188 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1438
timestamp 1681708930
transform 1 0 156 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1260
timestamp 1681708930
transform 1 0 156 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1234
timestamp 1681708930
transform 1 0 172 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_1439
timestamp 1681708930
transform 1 0 180 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1261
timestamp 1681708930
transform 1 0 180 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1202
timestamp 1681708930
transform 1 0 212 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_1368
timestamp 1681708930
transform 1 0 212 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1369
timestamp 1681708930
transform 1 0 220 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1235
timestamp 1681708930
transform 1 0 220 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_1440
timestamp 1681708930
transform 1 0 228 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1504
timestamp 1681708930
transform 1 0 212 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1505
timestamp 1681708930
transform 1 0 244 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1370
timestamp 1681708930
transform 1 0 276 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1441
timestamp 1681708930
transform 1 0 292 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1203
timestamp 1681708930
transform 1 0 300 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1204
timestamp 1681708930
transform 1 0 324 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_1353
timestamp 1681708930
transform 1 0 332 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1371
timestamp 1681708930
transform 1 0 300 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1372
timestamp 1681708930
transform 1 0 316 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1442
timestamp 1681708930
transform 1 0 308 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1443
timestamp 1681708930
transform 1 0 332 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1373
timestamp 1681708930
transform 1 0 348 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1288
timestamp 1681708930
transform 1 0 364 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1183
timestamp 1681708930
transform 1 0 380 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_1374
timestamp 1681708930
transform 1 0 380 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1444
timestamp 1681708930
transform 1 0 388 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1173
timestamp 1681708930
transform 1 0 444 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1184
timestamp 1681708930
transform 1 0 436 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1174
timestamp 1681708930
transform 1 0 492 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1185
timestamp 1681708930
transform 1 0 484 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1205
timestamp 1681708930
transform 1 0 444 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1206
timestamp 1681708930
transform 1 0 460 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_1375
timestamp 1681708930
transform 1 0 444 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1218
timestamp 1681708930
transform 1 0 468 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1236
timestamp 1681708930
transform 1 0 412 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1237
timestamp 1681708930
transform 1 0 444 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_1376
timestamp 1681708930
transform 1 0 484 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1445
timestamp 1681708930
transform 1 0 460 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1446
timestamp 1681708930
transform 1 0 476 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1262
timestamp 1681708930
transform 1 0 444 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1289
timestamp 1681708930
transform 1 0 436 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1238
timestamp 1681708930
transform 1 0 484 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1239
timestamp 1681708930
transform 1 0 500 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_1506
timestamp 1681708930
transform 1 0 476 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1507
timestamp 1681708930
transform 1 0 484 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_1290
timestamp 1681708930
transform 1 0 468 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1263
timestamp 1681708930
transform 1 0 492 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_1354
timestamp 1681708930
transform 1 0 516 0 1 1745
box -2 -2 2 2
use M3_M2  M3_M2_1219
timestamp 1681708930
transform 1 0 516 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_1377
timestamp 1681708930
transform 1 0 532 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1175
timestamp 1681708930
transform 1 0 548 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1186
timestamp 1681708930
transform 1 0 580 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_1355
timestamp 1681708930
transform 1 0 580 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1356
timestamp 1681708930
transform 1 0 588 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1378
timestamp 1681708930
transform 1 0 564 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1240
timestamp 1681708930
transform 1 0 540 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_1447
timestamp 1681708930
transform 1 0 548 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1241
timestamp 1681708930
transform 1 0 556 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1315
timestamp 1681708930
transform 1 0 564 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1187
timestamp 1681708930
transform 1 0 596 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1207
timestamp 1681708930
transform 1 0 612 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_1379
timestamp 1681708930
transform 1 0 612 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1220
timestamp 1681708930
transform 1 0 620 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1176
timestamp 1681708930
transform 1 0 652 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1188
timestamp 1681708930
transform 1 0 660 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1208
timestamp 1681708930
transform 1 0 644 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_1380
timestamp 1681708930
transform 1 0 628 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1381
timestamp 1681708930
transform 1 0 644 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1448
timestamp 1681708930
transform 1 0 612 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1242
timestamp 1681708930
transform 1 0 620 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1243
timestamp 1681708930
transform 1 0 636 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1264
timestamp 1681708930
transform 1 0 612 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1291
timestamp 1681708930
transform 1 0 604 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_1508
timestamp 1681708930
transform 1 0 636 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1528
timestamp 1681708930
transform 1 0 636 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_1316
timestamp 1681708930
transform 1 0 636 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1327
timestamp 1681708930
transform 1 0 628 0 1 1685
box -3 -3 3 3
use M2_M1  M2_M1_1509
timestamp 1681708930
transform 1 0 660 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_1265
timestamp 1681708930
transform 1 0 668 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1221
timestamp 1681708930
transform 1 0 684 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_1510
timestamp 1681708930
transform 1 0 676 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_1292
timestamp 1681708930
transform 1 0 660 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_1529
timestamp 1681708930
transform 1 0 668 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_1449
timestamp 1681708930
transform 1 0 692 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1293
timestamp 1681708930
transform 1 0 692 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1328
timestamp 1681708930
transform 1 0 708 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1294
timestamp 1681708930
transform 1 0 724 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1222
timestamp 1681708930
transform 1 0 740 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_1450
timestamp 1681708930
transform 1 0 740 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1317
timestamp 1681708930
transform 1 0 732 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1244
timestamp 1681708930
transform 1 0 748 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_1511
timestamp 1681708930
transform 1 0 748 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1451
timestamp 1681708930
transform 1 0 764 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1295
timestamp 1681708930
transform 1 0 764 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_1530
timestamp 1681708930
transform 1 0 772 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_1382
timestamp 1681708930
transform 1 0 852 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1383
timestamp 1681708930
transform 1 0 860 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1452
timestamp 1681708930
transform 1 0 860 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1266
timestamp 1681708930
transform 1 0 860 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_1384
timestamp 1681708930
transform 1 0 924 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1223
timestamp 1681708930
transform 1 0 940 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_1385
timestamp 1681708930
transform 1 0 948 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1453
timestamp 1681708930
transform 1 0 940 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1209
timestamp 1681708930
transform 1 0 996 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_1386
timestamp 1681708930
transform 1 0 996 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1387
timestamp 1681708930
transform 1 0 1004 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1454
timestamp 1681708930
transform 1 0 972 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1455
timestamp 1681708930
transform 1 0 980 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1267
timestamp 1681708930
transform 1 0 980 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1189
timestamp 1681708930
transform 1 0 1036 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1190
timestamp 1681708930
transform 1 0 1076 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1210
timestamp 1681708930
transform 1 0 1068 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_1388
timestamp 1681708930
transform 1 0 1036 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1389
timestamp 1681708930
transform 1 0 1052 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1390
timestamp 1681708930
transform 1 0 1060 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1456
timestamp 1681708930
transform 1 0 1044 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1245
timestamp 1681708930
transform 1 0 1052 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1268
timestamp 1681708930
transform 1 0 1044 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_1457
timestamp 1681708930
transform 1 0 1068 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1391
timestamp 1681708930
transform 1 0 1076 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1191
timestamp 1681708930
transform 1 0 1116 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_1392
timestamp 1681708930
transform 1 0 1108 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1393
timestamp 1681708930
transform 1 0 1116 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1458
timestamp 1681708930
transform 1 0 1100 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1246
timestamp 1681708930
transform 1 0 1108 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1224
timestamp 1681708930
transform 1 0 1124 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_1394
timestamp 1681708930
transform 1 0 1140 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1395
timestamp 1681708930
transform 1 0 1156 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1396
timestamp 1681708930
transform 1 0 1172 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1459
timestamp 1681708930
transform 1 0 1116 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1460
timestamp 1681708930
transform 1 0 1124 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1461
timestamp 1681708930
transform 1 0 1132 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1462
timestamp 1681708930
transform 1 0 1148 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1247
timestamp 1681708930
transform 1 0 1156 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_1463
timestamp 1681708930
transform 1 0 1164 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1296
timestamp 1681708930
transform 1 0 1164 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1297
timestamp 1681708930
transform 1 0 1180 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_1464
timestamp 1681708930
transform 1 0 1196 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1269
timestamp 1681708930
transform 1 0 1196 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1177
timestamp 1681708930
transform 1 0 1292 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1211
timestamp 1681708930
transform 1 0 1300 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_1397
timestamp 1681708930
transform 1 0 1212 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1225
timestamp 1681708930
transform 1 0 1236 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_1398
timestamp 1681708930
transform 1 0 1300 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1248
timestamp 1681708930
transform 1 0 1212 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_1465
timestamp 1681708930
transform 1 0 1236 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1466
timestamp 1681708930
transform 1 0 1292 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1270
timestamp 1681708930
transform 1 0 1236 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1298
timestamp 1681708930
transform 1 0 1244 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_1357
timestamp 1681708930
transform 1 0 1316 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1399
timestamp 1681708930
transform 1 0 1316 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1249
timestamp 1681708930
transform 1 0 1316 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_1467
timestamp 1681708930
transform 1 0 1324 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1212
timestamp 1681708930
transform 1 0 1420 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_1400
timestamp 1681708930
transform 1 0 1332 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1401
timestamp 1681708930
transform 1 0 1364 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1402
timestamp 1681708930
transform 1 0 1380 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1403
timestamp 1681708930
transform 1 0 1396 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1404
timestamp 1681708930
transform 1 0 1412 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1405
timestamp 1681708930
transform 1 0 1420 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1468
timestamp 1681708930
transform 1 0 1332 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1469
timestamp 1681708930
transform 1 0 1340 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1470
timestamp 1681708930
transform 1 0 1356 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1250
timestamp 1681708930
transform 1 0 1364 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1251
timestamp 1681708930
transform 1 0 1380 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_1471
timestamp 1681708930
transform 1 0 1388 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1299
timestamp 1681708930
transform 1 0 1332 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1226
timestamp 1681708930
transform 1 0 1444 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1252
timestamp 1681708930
transform 1 0 1452 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1192
timestamp 1681708930
transform 1 0 1524 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_1406
timestamp 1681708930
transform 1 0 1508 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1472
timestamp 1681708930
transform 1 0 1460 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1473
timestamp 1681708930
transform 1 0 1468 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1474
timestamp 1681708930
transform 1 0 1484 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1271
timestamp 1681708930
transform 1 0 1412 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1272
timestamp 1681708930
transform 1 0 1444 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_1512
timestamp 1681708930
transform 1 0 1452 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_1273
timestamp 1681708930
transform 1 0 1460 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_1513
timestamp 1681708930
transform 1 0 1476 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_1274
timestamp 1681708930
transform 1 0 1484 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1227
timestamp 1681708930
transform 1 0 1516 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_1475
timestamp 1681708930
transform 1 0 1516 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1514
timestamp 1681708930
transform 1 0 1500 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_1300
timestamp 1681708930
transform 1 0 1468 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_1531
timestamp 1681708930
transform 1 0 1484 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_1301
timestamp 1681708930
transform 1 0 1492 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1329
timestamp 1681708930
transform 1 0 1476 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1253
timestamp 1681708930
transform 1 0 1532 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_1515
timestamp 1681708930
transform 1 0 1532 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1407
timestamp 1681708930
transform 1 0 1548 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1330
timestamp 1681708930
transform 1 0 1556 0 1 1685
box -3 -3 3 3
use M2_M1  M2_M1_1408
timestamp 1681708930
transform 1 0 1588 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1331
timestamp 1681708930
transform 1 0 1588 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1193
timestamp 1681708930
transform 1 0 1604 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_1409
timestamp 1681708930
transform 1 0 1644 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1410
timestamp 1681708930
transform 1 0 1652 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1476
timestamp 1681708930
transform 1 0 1612 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1411
timestamp 1681708930
transform 1 0 1700 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1477
timestamp 1681708930
transform 1 0 1676 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1275
timestamp 1681708930
transform 1 0 1644 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1276
timestamp 1681708930
transform 1 0 1676 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1318
timestamp 1681708930
transform 1 0 1668 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1194
timestamp 1681708930
transform 1 0 1772 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_1412
timestamp 1681708930
transform 1 0 1756 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1478
timestamp 1681708930
transform 1 0 1732 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1479
timestamp 1681708930
transform 1 0 1740 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1254
timestamp 1681708930
transform 1 0 1756 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1195
timestamp 1681708930
transform 1 0 1844 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_1413
timestamp 1681708930
transform 1 0 1812 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1480
timestamp 1681708930
transform 1 0 1788 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1481
timestamp 1681708930
transform 1 0 1796 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1277
timestamp 1681708930
transform 1 0 1764 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1278
timestamp 1681708930
transform 1 0 1796 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1319
timestamp 1681708930
transform 1 0 1740 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_1414
timestamp 1681708930
transform 1 0 1868 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1415
timestamp 1681708930
transform 1 0 1876 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1482
timestamp 1681708930
transform 1 0 1844 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1255
timestamp 1681708930
transform 1 0 1876 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_1483
timestamp 1681708930
transform 1 0 1900 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1484
timestamp 1681708930
transform 1 0 1908 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1302
timestamp 1681708930
transform 1 0 1788 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1303
timestamp 1681708930
transform 1 0 1812 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1304
timestamp 1681708930
transform 1 0 1844 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1332
timestamp 1681708930
transform 1 0 1780 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1279
timestamp 1681708930
transform 1 0 1900 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1320
timestamp 1681708930
transform 1 0 1844 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1321
timestamp 1681708930
transform 1 0 1876 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_1416
timestamp 1681708930
transform 1 0 1932 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1485
timestamp 1681708930
transform 1 0 1964 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1178
timestamp 1681708930
transform 1 0 1996 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_1417
timestamp 1681708930
transform 1 0 1996 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1418
timestamp 1681708930
transform 1 0 2052 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1419
timestamp 1681708930
transform 1 0 2060 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1486
timestamp 1681708930
transform 1 0 2020 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1487
timestamp 1681708930
transform 1 0 2028 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1420
timestamp 1681708930
transform 1 0 2076 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1488
timestamp 1681708930
transform 1 0 2068 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1489
timestamp 1681708930
transform 1 0 2108 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1358
timestamp 1681708930
transform 1 0 2132 0 1 1745
box -2 -2 2 2
use M3_M2  M3_M2_1228
timestamp 1681708930
transform 1 0 2132 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_1421
timestamp 1681708930
transform 1 0 2148 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1490
timestamp 1681708930
transform 1 0 2132 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1256
timestamp 1681708930
transform 1 0 2164 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_1516
timestamp 1681708930
transform 1 0 2140 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_1305
timestamp 1681708930
transform 1 0 2116 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1280
timestamp 1681708930
transform 1 0 2148 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_1517
timestamp 1681708930
transform 1 0 2164 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1532
timestamp 1681708930
transform 1 0 2140 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_1306
timestamp 1681708930
transform 1 0 2164 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_1518
timestamp 1681708930
transform 1 0 2188 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_1229
timestamp 1681708930
transform 1 0 2220 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_1422
timestamp 1681708930
transform 1 0 2228 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1491
timestamp 1681708930
transform 1 0 2204 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1281
timestamp 1681708930
transform 1 0 2204 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_1519
timestamp 1681708930
transform 1 0 2220 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_1307
timestamp 1681708930
transform 1 0 2204 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_1533
timestamp 1681708930
transform 1 0 2212 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_1322
timestamp 1681708930
transform 1 0 2212 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1179
timestamp 1681708930
transform 1 0 2332 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1180
timestamp 1681708930
transform 1 0 2364 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1213
timestamp 1681708930
transform 1 0 2252 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1214
timestamp 1681708930
transform 1 0 2268 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1215
timestamp 1681708930
transform 1 0 2292 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_1492
timestamp 1681708930
transform 1 0 2236 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1493
timestamp 1681708930
transform 1 0 2244 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1282
timestamp 1681708930
transform 1 0 2236 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1323
timestamp 1681708930
transform 1 0 2244 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_1423
timestamp 1681708930
transform 1 0 2252 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1424
timestamp 1681708930
transform 1 0 2292 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1494
timestamp 1681708930
transform 1 0 2268 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1257
timestamp 1681708930
transform 1 0 2292 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1196
timestamp 1681708930
transform 1 0 2356 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1216
timestamp 1681708930
transform 1 0 2380 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1197
timestamp 1681708930
transform 1 0 2396 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_1359
timestamp 1681708930
transform 1 0 2388 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1425
timestamp 1681708930
transform 1 0 2340 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1426
timestamp 1681708930
transform 1 0 2356 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1427
timestamp 1681708930
transform 1 0 2380 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1428
timestamp 1681708930
transform 1 0 2388 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1495
timestamp 1681708930
transform 1 0 2316 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1496
timestamp 1681708930
transform 1 0 2324 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1520
timestamp 1681708930
transform 1 0 2260 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_1283
timestamp 1681708930
transform 1 0 2268 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_1521
timestamp 1681708930
transform 1 0 2284 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_1308
timestamp 1681708930
transform 1 0 2260 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_1534
timestamp 1681708930
transform 1 0 2276 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_1497
timestamp 1681708930
transform 1 0 2356 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_1309
timestamp 1681708930
transform 1 0 2340 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1310
timestamp 1681708930
transform 1 0 2364 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1333
timestamp 1681708930
transform 1 0 2324 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1334
timestamp 1681708930
transform 1 0 2356 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1198
timestamp 1681708930
transform 1 0 2436 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1230
timestamp 1681708930
transform 1 0 2428 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1199
timestamp 1681708930
transform 1 0 2492 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_1360
timestamp 1681708930
transform 1 0 2492 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1429
timestamp 1681708930
transform 1 0 2452 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1430
timestamp 1681708930
transform 1 0 2476 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1498
timestamp 1681708930
transform 1 0 2444 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1522
timestamp 1681708930
transform 1 0 2428 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_1311
timestamp 1681708930
transform 1 0 2428 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1258
timestamp 1681708930
transform 1 0 2452 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1231
timestamp 1681708930
transform 1 0 2492 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_1361
timestamp 1681708930
transform 1 0 2508 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1431
timestamp 1681708930
transform 1 0 2500 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1259
timestamp 1681708930
transform 1 0 2484 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_1523
timestamp 1681708930
transform 1 0 2460 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_1284
timestamp 1681708930
transform 1 0 2476 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_1499
timestamp 1681708930
transform 1 0 2508 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1524
timestamp 1681708930
transform 1 0 2484 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1535
timestamp 1681708930
transform 1 0 2468 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_1324
timestamp 1681708930
transform 1 0 2468 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1285
timestamp 1681708930
transform 1 0 2500 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1335
timestamp 1681708930
transform 1 0 2484 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1312
timestamp 1681708930
transform 1 0 2508 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_1362
timestamp 1681708930
transform 1 0 2524 0 1 1745
box -2 -2 2 2
use M3_M2  M3_M2_1336
timestamp 1681708930
transform 1 0 2516 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1232
timestamp 1681708930
transform 1 0 2532 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1217
timestamp 1681708930
transform 1 0 2572 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_1432
timestamp 1681708930
transform 1 0 2540 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1433
timestamp 1681708930
transform 1 0 2548 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1233
timestamp 1681708930
transform 1 0 2564 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_1434
timestamp 1681708930
transform 1 0 2572 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1500
timestamp 1681708930
transform 1 0 2532 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1501
timestamp 1681708930
transform 1 0 2540 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1435
timestamp 1681708930
transform 1 0 2596 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1502
timestamp 1681708930
transform 1 0 2588 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1525
timestamp 1681708930
transform 1 0 2572 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_1313
timestamp 1681708930
transform 1 0 2572 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_1526
timestamp 1681708930
transform 1 0 2604 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_1314
timestamp 1681708930
transform 1 0 2604 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1325
timestamp 1681708930
transform 1 0 2596 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1337
timestamp 1681708930
transform 1 0 2580 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1338
timestamp 1681708930
transform 1 0 2604 0 1 1685
box -3 -3 3 3
use M2_M1  M2_M1_1436
timestamp 1681708930
transform 1 0 2636 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1527
timestamp 1681708930
transform 1 0 2636 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1536
timestamp 1681708930
transform 1 0 2628 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_1326
timestamp 1681708930
transform 1 0 2636 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1339
timestamp 1681708930
transform 1 0 2644 0 1 1685
box -3 -3 3 3
use top_mod_new_VIA0  top_mod_new_VIA0_18
timestamp 1681708930
transform 1 0 24 0 1 1670
box -10 -3 10 3
use FILL  FILL_438
timestamp 1681708930
transform 1 0 72 0 -1 1770
box -8 -3 16 105
use FILL  FILL_440
timestamp 1681708930
transform 1 0 80 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_30
timestamp 1681708930
transform 1 0 88 0 -1 1770
box -8 -3 32 105
use FILL  FILL_445
timestamp 1681708930
transform 1 0 112 0 -1 1770
box -8 -3 16 105
use NAND2X1  NAND2X1_44
timestamp 1681708930
transform 1 0 120 0 -1 1770
box -8 -3 32 105
use FILL  FILL_450
timestamp 1681708930
transform 1 0 144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_451
timestamp 1681708930
transform 1 0 152 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_32
timestamp 1681708930
transform -1 0 184 0 -1 1770
box -8 -3 32 105
use OAI21X1  OAI21X1_41
timestamp 1681708930
transform 1 0 184 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_42
timestamp 1681708930
transform 1 0 216 0 -1 1770
box -8 -3 34 105
use FILL  FILL_452
timestamp 1681708930
transform 1 0 248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_453
timestamp 1681708930
transform 1 0 256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_454
timestamp 1681708930
transform 1 0 264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_455
timestamp 1681708930
transform 1 0 272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_456
timestamp 1681708930
transform 1 0 280 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_78
timestamp 1681708930
transform -1 0 304 0 -1 1770
box -9 -3 26 105
use AOI21X1  AOI21X1_17
timestamp 1681708930
transform 1 0 304 0 -1 1770
box -7 -3 39 105
use FILL  FILL_457
timestamp 1681708930
transform 1 0 336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_460
timestamp 1681708930
transform 1 0 344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_461
timestamp 1681708930
transform 1 0 352 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_33
timestamp 1681708930
transform 1 0 360 0 -1 1770
box -8 -3 32 105
use FILL  FILL_462
timestamp 1681708930
transform 1 0 384 0 -1 1770
box -8 -3 16 105
use XNOR2X1  XNOR2X1_16
timestamp 1681708930
transform 1 0 392 0 -1 1770
box -8 -3 64 105
use OAI21X1  OAI21X1_44
timestamp 1681708930
transform 1 0 448 0 -1 1770
box -8 -3 34 105
use NAND2X1  NAND2X1_46
timestamp 1681708930
transform -1 0 504 0 -1 1770
box -8 -3 32 105
use FILL  FILL_467
timestamp 1681708930
transform 1 0 504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_472
timestamp 1681708930
transform 1 0 512 0 -1 1770
box -8 -3 16 105
use FILL  FILL_473
timestamp 1681708930
transform 1 0 520 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_34
timestamp 1681708930
transform 1 0 528 0 -1 1770
box -8 -3 32 105
use AOI21X1  AOI21X1_20
timestamp 1681708930
transform 1 0 552 0 -1 1770
box -7 -3 39 105
use FILL  FILL_474
timestamp 1681708930
transform 1 0 584 0 -1 1770
box -8 -3 16 105
use FILL  FILL_475
timestamp 1681708930
transform 1 0 592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_476
timestamp 1681708930
transform 1 0 600 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_35
timestamp 1681708930
transform 1 0 608 0 -1 1770
box -8 -3 32 105
use NAND3X1  NAND3X1_42
timestamp 1681708930
transform 1 0 632 0 -1 1770
box -8 -3 40 105
use FILL  FILL_477
timestamp 1681708930
transform 1 0 664 0 -1 1770
box -8 -3 16 105
use FILL  FILL_478
timestamp 1681708930
transform 1 0 672 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_43
timestamp 1681708930
transform 1 0 680 0 -1 1770
box -8 -3 40 105
use FILL  FILL_479
timestamp 1681708930
transform 1 0 712 0 -1 1770
box -8 -3 16 105
use FILL  FILL_480
timestamp 1681708930
transform 1 0 720 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_81
timestamp 1681708930
transform 1 0 728 0 -1 1770
box -9 -3 26 105
use FILL  FILL_481
timestamp 1681708930
transform 1 0 744 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_44
timestamp 1681708930
transform 1 0 752 0 -1 1770
box -8 -3 40 105
use FILL  FILL_482
timestamp 1681708930
transform 1 0 784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_484
timestamp 1681708930
transform 1 0 792 0 -1 1770
box -8 -3 16 105
use XNOR2X1  XNOR2X1_19
timestamp 1681708930
transform 1 0 800 0 -1 1770
box -8 -3 64 105
use XNOR2X1  XNOR2X1_20
timestamp 1681708930
transform 1 0 856 0 -1 1770
box -8 -3 64 105
use FILL  FILL_491
timestamp 1681708930
transform 1 0 912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_502
timestamp 1681708930
transform 1 0 920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_503
timestamp 1681708930
transform 1 0 928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_504
timestamp 1681708930
transform 1 0 936 0 -1 1770
box -8 -3 16 105
use XOR2X1  XOR2X1_53
timestamp 1681708930
transform 1 0 944 0 -1 1770
box -8 -3 64 105
use FILL  FILL_505
timestamp 1681708930
transform 1 0 1000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_506
timestamp 1681708930
transform 1 0 1008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_507
timestamp 1681708930
transform 1 0 1016 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_14
timestamp 1681708930
transform 1 0 1024 0 -1 1770
box -8 -3 46 105
use FILL  FILL_508
timestamp 1681708930
transform 1 0 1064 0 -1 1770
box -8 -3 16 105
use FILL  FILL_509
timestamp 1681708930
transform 1 0 1072 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_15
timestamp 1681708930
transform 1 0 1080 0 -1 1770
box -8 -3 46 105
use FILL  FILL_510
timestamp 1681708930
transform 1 0 1120 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_16
timestamp 1681708930
transform 1 0 1128 0 -1 1770
box -8 -3 46 105
use INVX2  INVX2_85
timestamp 1681708930
transform 1 0 1168 0 -1 1770
box -9 -3 26 105
use FILL  FILL_519
timestamp 1681708930
transform 1 0 1184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_521
timestamp 1681708930
transform 1 0 1192 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_35
timestamp 1681708930
transform 1 0 1200 0 -1 1770
box -8 -3 104 105
use NOR2X1  NOR2X1_36
timestamp 1681708930
transform -1 0 1320 0 -1 1770
box -8 -3 32 105
use INVX2  INVX2_89
timestamp 1681708930
transform -1 0 1336 0 -1 1770
box -9 -3 26 105
use AOI22X1  AOI22X1_17
timestamp 1681708930
transform -1 0 1376 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_18
timestamp 1681708930
transform -1 0 1416 0 -1 1770
box -8 -3 46 105
use INVX2  INVX2_90
timestamp 1681708930
transform 1 0 1416 0 -1 1770
box -9 -3 26 105
use M3_M2  M3_M2_1340
timestamp 1681708930
transform 1 0 1460 0 1 1675
box -3 -3 3 3
use NAND2X1  NAND2X1_47
timestamp 1681708930
transform 1 0 1432 0 -1 1770
box -8 -3 32 105
use INVX2  INVX2_93
timestamp 1681708930
transform 1 0 1456 0 -1 1770
box -9 -3 26 105
use NAND3X1  NAND3X1_49
timestamp 1681708930
transform 1 0 1472 0 -1 1770
box -8 -3 40 105
use OAI21X1  OAI21X1_47
timestamp 1681708930
transform 1 0 1504 0 -1 1770
box -8 -3 34 105
use M3_M2  M3_M2_1341
timestamp 1681708930
transform 1 0 1548 0 1 1675
box -3 -3 3 3
use FILL  FILL_557
timestamp 1681708930
transform 1 0 1536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_558
timestamp 1681708930
transform 1 0 1544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_559
timestamp 1681708930
transform 1 0 1552 0 -1 1770
box -8 -3 16 105
use FILL  FILL_560
timestamp 1681708930
transform 1 0 1560 0 -1 1770
box -8 -3 16 105
use FILL  FILL_561
timestamp 1681708930
transform 1 0 1568 0 -1 1770
box -8 -3 16 105
use FILL  FILL_562
timestamp 1681708930
transform 1 0 1576 0 -1 1770
box -8 -3 16 105
use FILL  FILL_563
timestamp 1681708930
transform 1 0 1584 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_1342
timestamp 1681708930
transform 1 0 1636 0 1 1675
box -3 -3 3 3
use XOR2X1  XOR2X1_54
timestamp 1681708930
transform -1 0 1648 0 -1 1770
box -8 -3 64 105
use M3_M2  M3_M2_1343
timestamp 1681708930
transform 1 0 1708 0 1 1675
box -3 -3 3 3
use XOR2X1  XOR2X1_55
timestamp 1681708930
transform 1 0 1648 0 -1 1770
box -8 -3 64 105
use XOR2X1  XOR2X1_56
timestamp 1681708930
transform 1 0 1704 0 -1 1770
box -8 -3 64 105
use XOR2X1  XOR2X1_57
timestamp 1681708930
transform 1 0 1760 0 -1 1770
box -8 -3 64 105
use XOR2X1  XOR2X1_58
timestamp 1681708930
transform 1 0 1816 0 -1 1770
box -8 -3 64 105
use XOR2X1  XOR2X1_59
timestamp 1681708930
transform 1 0 1872 0 -1 1770
box -8 -3 64 105
use FILL  FILL_564
timestamp 1681708930
transform 1 0 1928 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_1344
timestamp 1681708930
transform 1 0 1964 0 1 1675
box -3 -3 3 3
use XOR2X1  XOR2X1_61
timestamp 1681708930
transform 1 0 1936 0 -1 1770
box -8 -3 64 105
use M3_M2  M3_M2_1345
timestamp 1681708930
transform 1 0 2004 0 1 1675
box -3 -3 3 3
use FILL  FILL_570
timestamp 1681708930
transform 1 0 1992 0 -1 1770
box -8 -3 16 105
use XOR2X1  XOR2X1_62
timestamp 1681708930
transform -1 0 2056 0 -1 1770
box -8 -3 64 105
use INVX2  INVX2_94
timestamp 1681708930
transform 1 0 2056 0 -1 1770
box -9 -3 26 105
use FILL  FILL_571
timestamp 1681708930
transform 1 0 2072 0 -1 1770
box -8 -3 16 105
use FILL  FILL_572
timestamp 1681708930
transform 1 0 2080 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_1346
timestamp 1681708930
transform 1 0 2100 0 1 1675
box -3 -3 3 3
use FILL  FILL_573
timestamp 1681708930
transform 1 0 2088 0 -1 1770
box -8 -3 16 105
use FILL  FILL_574
timestamp 1681708930
transform 1 0 2096 0 -1 1770
box -8 -3 16 105
use AOI21X1  AOI21X1_21
timestamp 1681708930
transform 1 0 2104 0 -1 1770
box -7 -3 39 105
use NAND3X1  NAND3X1_52
timestamp 1681708930
transform 1 0 2136 0 -1 1770
box -8 -3 40 105
use FILL  FILL_585
timestamp 1681708930
transform 1 0 2168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_586
timestamp 1681708930
transform 1 0 2176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_587
timestamp 1681708930
transform 1 0 2184 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_53
timestamp 1681708930
transform 1 0 2192 0 -1 1770
box -8 -3 40 105
use INVX2  INVX2_98
timestamp 1681708930
transform 1 0 2224 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_99
timestamp 1681708930
transform -1 0 2256 0 -1 1770
box -9 -3 26 105
use NAND3X1  NAND3X1_54
timestamp 1681708930
transform 1 0 2256 0 -1 1770
box -8 -3 40 105
use XOR2X1  XOR2X1_63
timestamp 1681708930
transform 1 0 2288 0 -1 1770
box -8 -3 64 105
use INVX2  INVX2_100
timestamp 1681708930
transform -1 0 2360 0 -1 1770
box -9 -3 26 105
use OR2X1  OR2X1_9
timestamp 1681708930
transform -1 0 2392 0 -1 1770
box -8 -3 40 105
use FILL  FILL_588
timestamp 1681708930
transform 1 0 2392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_589
timestamp 1681708930
transform 1 0 2400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_590
timestamp 1681708930
transform 1 0 2408 0 -1 1770
box -8 -3 16 105
use FILL  FILL_591
timestamp 1681708930
transform 1 0 2416 0 -1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_50
timestamp 1681708930
transform -1 0 2456 0 -1 1770
box -8 -3 34 105
use NAND3X1  NAND3X1_55
timestamp 1681708930
transform -1 0 2488 0 -1 1770
box -8 -3 40 105
use NOR2X1  NOR2X1_40
timestamp 1681708930
transform -1 0 2512 0 -1 1770
box -8 -3 32 105
use FILL  FILL_592
timestamp 1681708930
transform 1 0 2512 0 -1 1770
box -8 -3 16 105
use FILL  FILL_593
timestamp 1681708930
transform 1 0 2520 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_101
timestamp 1681708930
transform -1 0 2544 0 -1 1770
box -9 -3 26 105
use NOR2X1  NOR2X1_41
timestamp 1681708930
transform -1 0 2568 0 -1 1770
box -8 -3 32 105
use OAI21X1  OAI21X1_51
timestamp 1681708930
transform -1 0 2600 0 -1 1770
box -8 -3 34 105
use FILL  FILL_594
timestamp 1681708930
transform 1 0 2600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_595
timestamp 1681708930
transform 1 0 2608 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_56
timestamp 1681708930
transform -1 0 2648 0 -1 1770
box -8 -3 40 105
use FILL  FILL_596
timestamp 1681708930
transform 1 0 2648 0 -1 1770
box -8 -3 16 105
use FILL  FILL_598
timestamp 1681708930
transform 1 0 2656 0 -1 1770
box -8 -3 16 105
use top_mod_new_VIA0  top_mod_new_VIA0_19
timestamp 1681708930
transform 1 0 2712 0 1 1670
box -10 -3 10 3
use M2_M1  M2_M1_1565
timestamp 1681708930
transform 1 0 100 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1630
timestamp 1681708930
transform 1 0 108 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1537
timestamp 1681708930
transform 1 0 132 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_1547
timestamp 1681708930
transform 1 0 140 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1696
timestamp 1681708930
transform 1 0 148 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_1404
timestamp 1681708930
transform 1 0 164 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1566
timestamp 1681708930
transform 1 0 164 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1347
timestamp 1681708930
transform 1 0 188 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1363
timestamp 1681708930
transform 1 0 212 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_1538
timestamp 1681708930
transform 1 0 188 0 1 1635
box -2 -2 2 2
use M3_M2  M3_M2_1377
timestamp 1681708930
transform 1 0 196 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_1548
timestamp 1681708930
transform 1 0 196 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1567
timestamp 1681708930
transform 1 0 180 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1568
timestamp 1681708930
transform 1 0 204 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1364
timestamp 1681708930
transform 1 0 244 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1378
timestamp 1681708930
transform 1 0 244 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_1539
timestamp 1681708930
transform 1 0 252 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_1549
timestamp 1681708930
transform 1 0 236 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_1405
timestamp 1681708930
transform 1 0 252 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1569
timestamp 1681708930
transform 1 0 228 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1570
timestamp 1681708930
transform 1 0 244 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1631
timestamp 1681708930
transform 1 0 212 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1697
timestamp 1681708930
transform 1 0 228 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_1477
timestamp 1681708930
transform 1 0 236 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1379
timestamp 1681708930
transform 1 0 284 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_1540
timestamp 1681708930
transform 1 0 292 0 1 1635
box -2 -2 2 2
use M3_M2  M3_M2_1380
timestamp 1681708930
transform 1 0 300 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_1550
timestamp 1681708930
transform 1 0 268 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1551
timestamp 1681708930
transform 1 0 276 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_1470
timestamp 1681708930
transform 1 0 268 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1406
timestamp 1681708930
transform 1 0 284 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1541
timestamp 1681708930
transform 1 0 332 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_1552
timestamp 1681708930
transform 1 0 300 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1571
timestamp 1681708930
transform 1 0 284 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1407
timestamp 1681708930
transform 1 0 316 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1553
timestamp 1681708930
transform 1 0 324 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_1408
timestamp 1681708930
transform 1 0 332 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1441
timestamp 1681708930
transform 1 0 324 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1442
timestamp 1681708930
transform 1 0 340 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1632
timestamp 1681708930
transform 1 0 308 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1478
timestamp 1681708930
transform 1 0 308 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1498
timestamp 1681708930
transform 1 0 332 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1409
timestamp 1681708930
transform 1 0 356 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1633
timestamp 1681708930
transform 1 0 356 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1479
timestamp 1681708930
transform 1 0 356 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1499
timestamp 1681708930
transform 1 0 356 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_1554
timestamp 1681708930
transform 1 0 364 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_1443
timestamp 1681708930
transform 1 0 364 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1381
timestamp 1681708930
transform 1 0 388 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1410
timestamp 1681708930
transform 1 0 380 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1572
timestamp 1681708930
transform 1 0 380 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1573
timestamp 1681708930
transform 1 0 396 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1444
timestamp 1681708930
transform 1 0 404 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1634
timestamp 1681708930
transform 1 0 388 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1471
timestamp 1681708930
transform 1 0 396 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_1635
timestamp 1681708930
transform 1 0 404 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1500
timestamp 1681708930
transform 1 0 396 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1365
timestamp 1681708930
transform 1 0 428 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_1574
timestamp 1681708930
transform 1 0 420 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1382
timestamp 1681708930
transform 1 0 452 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_1575
timestamp 1681708930
transform 1 0 444 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1636
timestamp 1681708930
transform 1 0 428 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1480
timestamp 1681708930
transform 1 0 420 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1351
timestamp 1681708930
transform 1 0 484 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1411
timestamp 1681708930
transform 1 0 476 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1637
timestamp 1681708930
transform 1 0 468 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1638
timestamp 1681708930
transform 1 0 476 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1366
timestamp 1681708930
transform 1 0 524 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1445
timestamp 1681708930
transform 1 0 524 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1472
timestamp 1681708930
transform 1 0 492 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_1639
timestamp 1681708930
transform 1 0 540 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1481
timestamp 1681708930
transform 1 0 540 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1383
timestamp 1681708930
transform 1 0 556 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_1640
timestamp 1681708930
transform 1 0 556 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1367
timestamp 1681708930
transform 1 0 604 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_1576
timestamp 1681708930
transform 1 0 572 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1577
timestamp 1681708930
transform 1 0 580 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1578
timestamp 1681708930
transform 1 0 604 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1641
timestamp 1681708930
transform 1 0 588 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1482
timestamp 1681708930
transform 1 0 572 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1501
timestamp 1681708930
transform 1 0 588 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1384
timestamp 1681708930
transform 1 0 644 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1352
timestamp 1681708930
transform 1 0 684 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_1642
timestamp 1681708930
transform 1 0 644 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1643
timestamp 1681708930
transform 1 0 652 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1502
timestamp 1681708930
transform 1 0 652 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_1644
timestamp 1681708930
transform 1 0 700 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1483
timestamp 1681708930
transform 1 0 700 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1503
timestamp 1681708930
transform 1 0 708 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_1579
timestamp 1681708930
transform 1 0 724 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1473
timestamp 1681708930
transform 1 0 724 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1353
timestamp 1681708930
transform 1 0 828 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1385
timestamp 1681708930
transform 1 0 740 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1386
timestamp 1681708930
transform 1 0 756 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1412
timestamp 1681708930
transform 1 0 740 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1413
timestamp 1681708930
transform 1 0 780 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1580
timestamp 1681708930
transform 1 0 740 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1446
timestamp 1681708930
transform 1 0 756 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1581
timestamp 1681708930
transform 1 0 780 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1447
timestamp 1681708930
transform 1 0 804 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1582
timestamp 1681708930
transform 1 0 836 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1645
timestamp 1681708930
transform 1 0 732 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1448
timestamp 1681708930
transform 1 0 852 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1583
timestamp 1681708930
transform 1 0 860 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1449
timestamp 1681708930
transform 1 0 868 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1584
timestamp 1681708930
transform 1 0 884 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1646
timestamp 1681708930
transform 1 0 756 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1647
timestamp 1681708930
transform 1 0 844 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1648
timestamp 1681708930
transform 1 0 852 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1649
timestamp 1681708930
transform 1 0 868 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1650
timestamp 1681708930
transform 1 0 876 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1484
timestamp 1681708930
transform 1 0 844 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1504
timestamp 1681708930
transform 1 0 756 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1505
timestamp 1681708930
transform 1 0 836 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1348
timestamp 1681708930
transform 1 0 956 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1354
timestamp 1681708930
transform 1 0 908 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1355
timestamp 1681708930
transform 1 0 924 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1356
timestamp 1681708930
transform 1 0 940 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1387
timestamp 1681708930
transform 1 0 908 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1388
timestamp 1681708930
transform 1 0 932 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1414
timestamp 1681708930
transform 1 0 892 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1415
timestamp 1681708930
transform 1 0 932 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1416
timestamp 1681708930
transform 1 0 1028 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1585
timestamp 1681708930
transform 1 0 892 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1586
timestamp 1681708930
transform 1 0 932 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1587
timestamp 1681708930
transform 1 0 988 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1588
timestamp 1681708930
transform 1 0 1012 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1589
timestamp 1681708930
transform 1 0 1028 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1590
timestamp 1681708930
transform 1 0 1036 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1651
timestamp 1681708930
transform 1 0 908 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1474
timestamp 1681708930
transform 1 0 988 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_1652
timestamp 1681708930
transform 1 0 996 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1653
timestamp 1681708930
transform 1 0 1004 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1654
timestamp 1681708930
transform 1 0 1028 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1485
timestamp 1681708930
transform 1 0 884 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1486
timestamp 1681708930
transform 1 0 908 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1487
timestamp 1681708930
transform 1 0 980 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1488
timestamp 1681708930
transform 1 0 1028 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1450
timestamp 1681708930
transform 1 0 1052 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1655
timestamp 1681708930
transform 1 0 1044 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1389
timestamp 1681708930
transform 1 0 1108 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_1591
timestamp 1681708930
transform 1 0 1108 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1656
timestamp 1681708930
transform 1 0 1108 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1489
timestamp 1681708930
transform 1 0 1108 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1417
timestamp 1681708930
transform 1 0 1124 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1592
timestamp 1681708930
transform 1 0 1148 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1593
timestamp 1681708930
transform 1 0 1164 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1657
timestamp 1681708930
transform 1 0 1140 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1451
timestamp 1681708930
transform 1 0 1172 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1658
timestamp 1681708930
transform 1 0 1172 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1418
timestamp 1681708930
transform 1 0 1188 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1594
timestamp 1681708930
transform 1 0 1188 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1506
timestamp 1681708930
transform 1 0 1188 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1390
timestamp 1681708930
transform 1 0 1204 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_1659
timestamp 1681708930
transform 1 0 1204 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1391
timestamp 1681708930
transform 1 0 1292 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1419
timestamp 1681708930
transform 1 0 1268 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1452
timestamp 1681708930
transform 1 0 1260 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1420
timestamp 1681708930
transform 1 0 1300 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1421
timestamp 1681708930
transform 1 0 1316 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1595
timestamp 1681708930
transform 1 0 1268 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1596
timestamp 1681708930
transform 1 0 1284 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1453
timestamp 1681708930
transform 1 0 1292 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1597
timestamp 1681708930
transform 1 0 1300 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1660
timestamp 1681708930
transform 1 0 1252 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1661
timestamp 1681708930
transform 1 0 1260 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1662
timestamp 1681708930
transform 1 0 1276 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1663
timestamp 1681708930
transform 1 0 1300 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1664
timestamp 1681708930
transform 1 0 1316 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1490
timestamp 1681708930
transform 1 0 1300 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_1555
timestamp 1681708930
transform 1 0 1340 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_1454
timestamp 1681708930
transform 1 0 1340 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1368
timestamp 1681708930
transform 1 0 1356 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1491
timestamp 1681708930
transform 1 0 1348 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_1598
timestamp 1681708930
transform 1 0 1372 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1599
timestamp 1681708930
transform 1 0 1380 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1392
timestamp 1681708930
transform 1 0 1412 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_1665
timestamp 1681708930
transform 1 0 1404 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1422
timestamp 1681708930
transform 1 0 1420 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1556
timestamp 1681708930
transform 1 0 1428 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_1455
timestamp 1681708930
transform 1 0 1420 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1600
timestamp 1681708930
transform 1 0 1428 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1456
timestamp 1681708930
transform 1 0 1436 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1601
timestamp 1681708930
transform 1 0 1444 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1542
timestamp 1681708930
transform 1 0 1452 0 1 1635
box -2 -2 2 2
use M3_M2  M3_M2_1423
timestamp 1681708930
transform 1 0 1452 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1666
timestamp 1681708930
transform 1 0 1452 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1357
timestamp 1681708930
transform 1 0 1468 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1349
timestamp 1681708930
transform 1 0 1500 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1424
timestamp 1681708930
transform 1 0 1492 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1602
timestamp 1681708930
transform 1 0 1484 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1603
timestamp 1681708930
transform 1 0 1492 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1475
timestamp 1681708930
transform 1 0 1484 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1492
timestamp 1681708930
transform 1 0 1492 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1393
timestamp 1681708930
transform 1 0 1508 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1369
timestamp 1681708930
transform 1 0 1524 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_1543
timestamp 1681708930
transform 1 0 1524 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_1557
timestamp 1681708930
transform 1 0 1516 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_1425
timestamp 1681708930
transform 1 0 1524 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1457
timestamp 1681708930
transform 1 0 1516 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1667
timestamp 1681708930
transform 1 0 1508 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1507
timestamp 1681708930
transform 1 0 1500 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_1698
timestamp 1681708930
transform 1 0 1516 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_1350
timestamp 1681708930
transform 1 0 1580 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1358
timestamp 1681708930
transform 1 0 1556 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1394
timestamp 1681708930
transform 1 0 1548 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1370
timestamp 1681708930
transform 1 0 1596 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_1558
timestamp 1681708930
transform 1 0 1556 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_1371
timestamp 1681708930
transform 1 0 1652 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1372
timestamp 1681708930
transform 1 0 1700 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1395
timestamp 1681708930
transform 1 0 1676 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1426
timestamp 1681708930
transform 1 0 1620 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1427
timestamp 1681708930
transform 1 0 1652 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1604
timestamp 1681708930
transform 1 0 1540 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1458
timestamp 1681708930
transform 1 0 1556 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1605
timestamp 1681708930
transform 1 0 1564 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1459
timestamp 1681708930
transform 1 0 1588 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1606
timestamp 1681708930
transform 1 0 1620 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1668
timestamp 1681708930
transform 1 0 1564 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1493
timestamp 1681708930
transform 1 0 1564 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1508
timestamp 1681708930
transform 1 0 1540 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1460
timestamp 1681708930
transform 1 0 1636 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1607
timestamp 1681708930
transform 1 0 1676 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1669
timestamp 1681708930
transform 1 0 1612 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1670
timestamp 1681708930
transform 1 0 1620 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1509
timestamp 1681708930
transform 1 0 1596 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_1671
timestamp 1681708930
transform 1 0 1668 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1672
timestamp 1681708930
transform 1 0 1676 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1494
timestamp 1681708930
transform 1 0 1668 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1510
timestamp 1681708930
transform 1 0 1636 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1511
timestamp 1681708930
transform 1 0 1652 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1512
timestamp 1681708930
transform 1 0 1676 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1428
timestamp 1681708930
transform 1 0 1732 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1429
timestamp 1681708930
transform 1 0 1764 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1396
timestamp 1681708930
transform 1 0 1812 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1397
timestamp 1681708930
transform 1 0 1836 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_1608
timestamp 1681708930
transform 1 0 1764 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1673
timestamp 1681708930
transform 1 0 1732 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1513
timestamp 1681708930
transform 1 0 1724 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1461
timestamp 1681708930
transform 1 0 1780 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1609
timestamp 1681708930
transform 1 0 1812 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1610
timestamp 1681708930
transform 1 0 1820 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1674
timestamp 1681708930
transform 1 0 1780 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1675
timestamp 1681708930
transform 1 0 1788 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1373
timestamp 1681708930
transform 1 0 1900 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1398
timestamp 1681708930
transform 1 0 1892 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1430
timestamp 1681708930
transform 1 0 1868 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1611
timestamp 1681708930
transform 1 0 1868 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1462
timestamp 1681708930
transform 1 0 1876 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1676
timestamp 1681708930
transform 1 0 1836 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1514
timestamp 1681708930
transform 1 0 1876 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1359
timestamp 1681708930
transform 1 0 1924 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1360
timestamp 1681708930
transform 1 0 1972 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1361
timestamp 1681708930
transform 1 0 1988 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1362
timestamp 1681708930
transform 1 0 2004 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_1677
timestamp 1681708930
transform 1 0 1916 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1495
timestamp 1681708930
transform 1 0 1916 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1399
timestamp 1681708930
transform 1 0 2012 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_1612
timestamp 1681708930
transform 1 0 1956 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1613
timestamp 1681708930
transform 1 0 2012 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1614
timestamp 1681708930
transform 1 0 2020 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1678
timestamp 1681708930
transform 1 0 1932 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1496
timestamp 1681708930
transform 1 0 1980 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1515
timestamp 1681708930
transform 1 0 1924 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1516
timestamp 1681708930
transform 1 0 1956 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_1679
timestamp 1681708930
transform 1 0 2020 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1497
timestamp 1681708930
transform 1 0 2020 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1431
timestamp 1681708930
transform 1 0 2060 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1615
timestamp 1681708930
transform 1 0 2036 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1616
timestamp 1681708930
transform 1 0 2060 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1374
timestamp 1681708930
transform 1 0 2092 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1432
timestamp 1681708930
transform 1 0 2108 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1433
timestamp 1681708930
transform 1 0 2140 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1617
timestamp 1681708930
transform 1 0 2140 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1680
timestamp 1681708930
transform 1 0 2108 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1681
timestamp 1681708930
transform 1 0 2116 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1517
timestamp 1681708930
transform 1 0 2156 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1434
timestamp 1681708930
transform 1 0 2172 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1682
timestamp 1681708930
transform 1 0 2172 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1683
timestamp 1681708930
transform 1 0 2180 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1435
timestamp 1681708930
transform 1 0 2228 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1618
timestamp 1681708930
transform 1 0 2228 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1684
timestamp 1681708930
transform 1 0 2204 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1518
timestamp 1681708930
transform 1 0 2196 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1436
timestamp 1681708930
transform 1 0 2260 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1619
timestamp 1681708930
transform 1 0 2268 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1463
timestamp 1681708930
transform 1 0 2276 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1437
timestamp 1681708930
transform 1 0 2316 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1620
timestamp 1681708930
transform 1 0 2284 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1685
timestamp 1681708930
transform 1 0 2276 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1686
timestamp 1681708930
transform 1 0 2284 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1519
timestamp 1681708930
transform 1 0 2268 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_1621
timestamp 1681708930
transform 1 0 2332 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1520
timestamp 1681708930
transform 1 0 2308 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_1544
timestamp 1681708930
transform 1 0 2356 0 1 1635
box -2 -2 2 2
use M3_M2  M3_M2_1400
timestamp 1681708930
transform 1 0 2364 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_1559
timestamp 1681708930
transform 1 0 2348 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1687
timestamp 1681708930
transform 1 0 2340 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1545
timestamp 1681708930
transform 1 0 2396 0 1 1635
box -2 -2 2 2
use M3_M2  M3_M2_1401
timestamp 1681708930
transform 1 0 2404 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_1560
timestamp 1681708930
transform 1 0 2372 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1561
timestamp 1681708930
transform 1 0 2380 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_1438
timestamp 1681708930
transform 1 0 2396 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_1562
timestamp 1681708930
transform 1 0 2404 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1622
timestamp 1681708930
transform 1 0 2364 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1464
timestamp 1681708930
transform 1 0 2380 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1623
timestamp 1681708930
transform 1 0 2396 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1476
timestamp 1681708930
transform 1 0 2372 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1465
timestamp 1681708930
transform 1 0 2404 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1563
timestamp 1681708930
transform 1 0 2436 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1546
timestamp 1681708930
transform 1 0 2452 0 1 1635
box -2 -2 2 2
use M3_M2  M3_M2_1402
timestamp 1681708930
transform 1 0 2468 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_1564
timestamp 1681708930
transform 1 0 2468 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_1439
timestamp 1681708930
transform 1 0 2476 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1466
timestamp 1681708930
transform 1 0 2452 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1624
timestamp 1681708930
transform 1 0 2460 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1625
timestamp 1681708930
transform 1 0 2476 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1375
timestamp 1681708930
transform 1 0 2516 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_1626
timestamp 1681708930
transform 1 0 2500 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1403
timestamp 1681708930
transform 1 0 2524 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_1627
timestamp 1681708930
transform 1 0 2524 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1376
timestamp 1681708930
transform 1 0 2548 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1440
timestamp 1681708930
transform 1 0 2588 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1467
timestamp 1681708930
transform 1 0 2548 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1468
timestamp 1681708930
transform 1 0 2580 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1628
timestamp 1681708930
transform 1 0 2588 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_1469
timestamp 1681708930
transform 1 0 2612 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_1629
timestamp 1681708930
transform 1 0 2636 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1688
timestamp 1681708930
transform 1 0 2500 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1689
timestamp 1681708930
transform 1 0 2508 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1690
timestamp 1681708930
transform 1 0 2532 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1691
timestamp 1681708930
transform 1 0 2540 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1692
timestamp 1681708930
transform 1 0 2548 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1699
timestamp 1681708930
transform 1 0 2524 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_1521
timestamp 1681708930
transform 1 0 2516 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_1700
timestamp 1681708930
transform 1 0 2548 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_1522
timestamp 1681708930
transform 1 0 2540 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_1693
timestamp 1681708930
transform 1 0 2604 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1694
timestamp 1681708930
transform 1 0 2612 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1695
timestamp 1681708930
transform 1 0 2668 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_1523
timestamp 1681708930
transform 1 0 2564 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1524
timestamp 1681708930
transform 1 0 2596 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1525
timestamp 1681708930
transform 1 0 2660 0 1 1585
box -3 -3 3 3
use top_mod_new_VIA0  top_mod_new_VIA0_20
timestamp 1681708930
transform 1 0 48 0 1 1570
box -10 -3 10 3
use FILL  FILL_599
timestamp 1681708930
transform 1 0 72 0 1 1570
box -8 -3 16 105
use FILL  FILL_600
timestamp 1681708930
transform 1 0 80 0 1 1570
box -8 -3 16 105
use FILL  FILL_601
timestamp 1681708930
transform 1 0 88 0 1 1570
box -8 -3 16 105
use AOI21X1  AOI21X1_25
timestamp 1681708930
transform 1 0 96 0 1 1570
box -7 -3 39 105
use FILL  FILL_602
timestamp 1681708930
transform 1 0 128 0 1 1570
box -8 -3 16 105
use FILL  FILL_603
timestamp 1681708930
transform 1 0 136 0 1 1570
box -8 -3 16 105
use FILL  FILL_604
timestamp 1681708930
transform 1 0 144 0 1 1570
box -8 -3 16 105
use FILL  FILL_605
timestamp 1681708930
transform 1 0 152 0 1 1570
box -8 -3 16 105
use FILL  FILL_606
timestamp 1681708930
transform 1 0 160 0 1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_57
timestamp 1681708930
transform 1 0 168 0 1 1570
box -8 -3 40 105
use AOI21X1  AOI21X1_26
timestamp 1681708930
transform 1 0 200 0 1 1570
box -7 -3 39 105
use NAND3X1  NAND3X1_58
timestamp 1681708930
transform 1 0 232 0 1 1570
box -8 -3 40 105
use FILL  FILL_607
timestamp 1681708930
transform 1 0 264 0 1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_59
timestamp 1681708930
transform 1 0 272 0 1 1570
box -8 -3 40 105
use INVX2  INVX2_102
timestamp 1681708930
transform 1 0 304 0 1 1570
box -9 -3 26 105
use M3_M2  M3_M2_1526
timestamp 1681708930
transform 1 0 348 0 1 1575
box -3 -3 3 3
use NAND3X1  NAND3X1_60
timestamp 1681708930
transform 1 0 320 0 1 1570
box -8 -3 40 105
use FILL  FILL_608
timestamp 1681708930
transform 1 0 352 0 1 1570
box -8 -3 16 105
use FILL  FILL_609
timestamp 1681708930
transform 1 0 360 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_103
timestamp 1681708930
transform 1 0 368 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_104
timestamp 1681708930
transform 1 0 384 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_105
timestamp 1681708930
transform 1 0 400 0 1 1570
box -9 -3 26 105
use FILL  FILL_610
timestamp 1681708930
transform 1 0 416 0 1 1570
box -8 -3 16 105
use BUFX2  BUFX2_1
timestamp 1681708930
transform -1 0 448 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_2
timestamp 1681708930
transform 1 0 448 0 1 1570
box -5 -3 28 105
use FILL  FILL_611
timestamp 1681708930
transform 1 0 472 0 1 1570
box -8 -3 16 105
use FILL  FILL_612
timestamp 1681708930
transform 1 0 480 0 1 1570
box -8 -3 16 105
use XNOR2X1  XNOR2X1_23
timestamp 1681708930
transform 1 0 488 0 1 1570
box -8 -3 64 105
use FILL  FILL_613
timestamp 1681708930
transform 1 0 544 0 1 1570
box -8 -3 16 105
use FILL  FILL_614
timestamp 1681708930
transform 1 0 552 0 1 1570
box -8 -3 16 105
use FILL  FILL_615
timestamp 1681708930
transform 1 0 560 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_1527
timestamp 1681708930
transform 1 0 604 0 1 1575
box -3 -3 3 3
use INVX2  INVX2_106
timestamp 1681708930
transform 1 0 568 0 1 1570
box -9 -3 26 105
use XNOR2X1  XNOR2X1_25
timestamp 1681708930
transform -1 0 640 0 1 1570
box -8 -3 64 105
use FILL  FILL_616
timestamp 1681708930
transform 1 0 640 0 1 1570
box -8 -3 16 105
use XOR2X1  XOR2X1_64
timestamp 1681708930
transform 1 0 648 0 1 1570
box -8 -3 64 105
use FILL  FILL_617
timestamp 1681708930
transform 1 0 704 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_1528
timestamp 1681708930
transform 1 0 724 0 1 1575
box -3 -3 3 3
use FILL  FILL_618
timestamp 1681708930
transform 1 0 712 0 1 1570
box -8 -3 16 105
use FILL  FILL_619
timestamp 1681708930
transform 1 0 720 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_1529
timestamp 1681708930
transform 1 0 748 0 1 1575
box -3 -3 3 3
use INVX2  INVX2_107
timestamp 1681708930
transform 1 0 728 0 1 1570
box -9 -3 26 105
use M3_M2  M3_M2_1530
timestamp 1681708930
transform 1 0 812 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_39
timestamp 1681708930
transform 1 0 744 0 1 1570
box -8 -3 104 105
use AOI22X1  AOI22X1_23
timestamp 1681708930
transform 1 0 840 0 1 1570
box -8 -3 46 105
use INVX2  INVX2_108
timestamp 1681708930
transform 1 0 880 0 1 1570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_40
timestamp 1681708930
transform 1 0 896 0 1 1570
box -8 -3 104 105
use M3_M2  M3_M2_1531
timestamp 1681708930
transform 1 0 1020 0 1 1575
box -3 -3 3 3
use AOI22X1  AOI22X1_24
timestamp 1681708930
transform 1 0 992 0 1 1570
box -8 -3 46 105
use M3_M2  M3_M2_1532
timestamp 1681708930
transform 1 0 1044 0 1 1575
box -3 -3 3 3
use FILL  FILL_620
timestamp 1681708930
transform 1 0 1032 0 1 1570
box -8 -3 16 105
use FILL  FILL_624
timestamp 1681708930
transform 1 0 1040 0 1 1570
box -8 -3 16 105
use FILL  FILL_625
timestamp 1681708930
transform 1 0 1048 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_1533
timestamp 1681708930
transform 1 0 1100 0 1 1575
box -3 -3 3 3
use XOR2X1  XOR2X1_67
timestamp 1681708930
transform -1 0 1112 0 1 1570
box -8 -3 64 105
use FILL  FILL_626
timestamp 1681708930
transform 1 0 1112 0 1 1570
box -8 -3 16 105
use FILL  FILL_627
timestamp 1681708930
transform 1 0 1120 0 1 1570
box -8 -3 16 105
use FILL  FILL_628
timestamp 1681708930
transform 1 0 1128 0 1 1570
box -8 -3 16 105
use FILL  FILL_629
timestamp 1681708930
transform 1 0 1136 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_28
timestamp 1681708930
transform 1 0 1144 0 1 1570
box -8 -3 46 105
use FILL  FILL_630
timestamp 1681708930
transform 1 0 1184 0 1 1570
box -8 -3 16 105
use FILL  FILL_631
timestamp 1681708930
transform 1 0 1192 0 1 1570
box -8 -3 16 105
use XOR2X1  XOR2X1_68
timestamp 1681708930
transform -1 0 1256 0 1 1570
box -8 -3 64 105
use OAI22X1  OAI22X1_20
timestamp 1681708930
transform 1 0 1256 0 1 1570
box -8 -3 46 105
use FILL  FILL_632
timestamp 1681708930
transform 1 0 1296 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_111
timestamp 1681708930
transform -1 0 1320 0 1 1570
box -9 -3 26 105
use NAND2X1  NAND2X1_48
timestamp 1681708930
transform 1 0 1320 0 1 1570
box -8 -3 32 105
use FILL  FILL_633
timestamp 1681708930
transform 1 0 1344 0 1 1570
box -8 -3 16 105
use FILL  FILL_634
timestamp 1681708930
transform 1 0 1352 0 1 1570
box -8 -3 16 105
use FILL  FILL_635
timestamp 1681708930
transform 1 0 1360 0 1 1570
box -8 -3 16 105
use FILL  FILL_636
timestamp 1681708930
transform 1 0 1368 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_112
timestamp 1681708930
transform -1 0 1392 0 1 1570
box -9 -3 26 105
use FILL  FILL_637
timestamp 1681708930
transform 1 0 1392 0 1 1570
box -8 -3 16 105
use FILL  FILL_638
timestamp 1681708930
transform 1 0 1400 0 1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_64
timestamp 1681708930
transform -1 0 1440 0 1 1570
box -8 -3 40 105
use FILL  FILL_639
timestamp 1681708930
transform 1 0 1440 0 1 1570
box -8 -3 16 105
use FILL  FILL_640
timestamp 1681708930
transform 1 0 1448 0 1 1570
box -8 -3 16 105
use AOI21X1  AOI21X1_27
timestamp 1681708930
transform 1 0 1456 0 1 1570
box -7 -3 39 105
use NOR2X1  NOR2X1_42
timestamp 1681708930
transform -1 0 1512 0 1 1570
box -8 -3 32 105
use FILL  FILL_641
timestamp 1681708930
transform 1 0 1512 0 1 1570
box -8 -3 16 105
use FILL  FILL_642
timestamp 1681708930
transform 1 0 1520 0 1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_65
timestamp 1681708930
transform 1 0 1528 0 1 1570
box -8 -3 40 105
use XNOR2X1  XNOR2X1_28
timestamp 1681708930
transform -1 0 1616 0 1 1570
box -8 -3 64 105
use XOR2X1  XOR2X1_69
timestamp 1681708930
transform -1 0 1672 0 1 1570
box -8 -3 64 105
use XOR2X1  XOR2X1_70
timestamp 1681708930
transform -1 0 1728 0 1 1570
box -8 -3 64 105
use XOR2X1  XOR2X1_71
timestamp 1681708930
transform 1 0 1728 0 1 1570
box -8 -3 64 105
use XOR2X1  XOR2X1_72
timestamp 1681708930
transform 1 0 1784 0 1 1570
box -8 -3 64 105
use XOR2X1  XOR2X1_73
timestamp 1681708930
transform 1 0 1840 0 1 1570
box -8 -3 64 105
use FILL  FILL_643
timestamp 1681708930
transform 1 0 1896 0 1 1570
box -8 -3 16 105
use FILL  FILL_650
timestamp 1681708930
transform 1 0 1904 0 1 1570
box -8 -3 16 105
use FILL  FILL_652
timestamp 1681708930
transform 1 0 1912 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_1534
timestamp 1681708930
transform 1 0 1940 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1535
timestamp 1681708930
transform 1 0 1964 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_43
timestamp 1681708930
transform 1 0 1920 0 1 1570
box -8 -3 104 105
use FILL  FILL_653
timestamp 1681708930
transform 1 0 2016 0 1 1570
box -8 -3 16 105
use FILL  FILL_654
timestamp 1681708930
transform 1 0 2024 0 1 1570
box -8 -3 16 105
use XOR2X1  XOR2X1_80
timestamp 1681708930
transform -1 0 2088 0 1 1570
box -8 -3 64 105
use FILL  FILL_655
timestamp 1681708930
transform 1 0 2088 0 1 1570
box -8 -3 16 105
use FILL  FILL_656
timestamp 1681708930
transform 1 0 2096 0 1 1570
box -8 -3 16 105
use FILL  FILL_657
timestamp 1681708930
transform 1 0 2104 0 1 1570
box -8 -3 16 105
use XOR2X1  XOR2X1_81
timestamp 1681708930
transform 1 0 2112 0 1 1570
box -8 -3 64 105
use FILL  FILL_658
timestamp 1681708930
transform 1 0 2168 0 1 1570
box -8 -3 16 105
use FILL  FILL_669
timestamp 1681708930
transform 1 0 2176 0 1 1570
box -8 -3 16 105
use FILL  FILL_670
timestamp 1681708930
transform 1 0 2184 0 1 1570
box -8 -3 16 105
use FILL  FILL_671
timestamp 1681708930
transform 1 0 2192 0 1 1570
box -8 -3 16 105
use XOR2X1  XOR2X1_83
timestamp 1681708930
transform 1 0 2200 0 1 1570
box -8 -3 64 105
use FILL  FILL_672
timestamp 1681708930
transform 1 0 2256 0 1 1570
box -8 -3 16 105
use FILL  FILL_673
timestamp 1681708930
transform 1 0 2264 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_1536
timestamp 1681708930
transform 1 0 2284 0 1 1575
box -3 -3 3 3
use FILL  FILL_674
timestamp 1681708930
transform 1 0 2272 0 1 1570
box -8 -3 16 105
use XOR2X1  XOR2X1_84
timestamp 1681708930
transform 1 0 2280 0 1 1570
box -8 -3 64 105
use FILL  FILL_675
timestamp 1681708930
transform 1 0 2336 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_1537
timestamp 1681708930
transform 1 0 2364 0 1 1575
box -3 -3 3 3
use NAND3X1  NAND3X1_67
timestamp 1681708930
transform -1 0 2376 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_68
timestamp 1681708930
transform -1 0 2408 0 1 1570
box -8 -3 40 105
use FILL  FILL_676
timestamp 1681708930
transform 1 0 2408 0 1 1570
box -8 -3 16 105
use FILL  FILL_677
timestamp 1681708930
transform 1 0 2416 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_1538
timestamp 1681708930
transform 1 0 2436 0 1 1575
box -3 -3 3 3
use FILL  FILL_678
timestamp 1681708930
transform 1 0 2424 0 1 1570
box -8 -3 16 105
use FILL  FILL_679
timestamp 1681708930
transform 1 0 2432 0 1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_69
timestamp 1681708930
transform -1 0 2472 0 1 1570
box -8 -3 40 105
use INVX2  INVX2_118
timestamp 1681708930
transform -1 0 2488 0 1 1570
box -9 -3 26 105
use FILL  FILL_680
timestamp 1681708930
transform 1 0 2488 0 1 1570
box -8 -3 16 105
use AOI21X1  AOI21X1_28
timestamp 1681708930
transform 1 0 2496 0 1 1570
box -7 -3 39 105
use M3_M2  M3_M2_1539
timestamp 1681708930
transform 1 0 2548 0 1 1575
box -3 -3 3 3
use NOR2X1  NOR2X1_44
timestamp 1681708930
transform -1 0 2552 0 1 1570
box -8 -3 32 105
use M3_M2  M3_M2_1540
timestamp 1681708930
transform 1 0 2604 0 1 1575
box -3 -3 3 3
use XNOR2X1  XNOR2X1_32
timestamp 1681708930
transform 1 0 2552 0 1 1570
box -8 -3 64 105
use XOR2X1  XOR2X1_85
timestamp 1681708930
transform -1 0 2664 0 1 1570
box -8 -3 64 105
use top_mod_new_VIA0  top_mod_new_VIA0_21
timestamp 1681708930
transform 1 0 2688 0 1 1570
box -10 -3 10 3
use M3_M2  M3_M2_1591
timestamp 1681708930
transform 1 0 84 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1704
timestamp 1681708930
transform 1 0 84 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_1592
timestamp 1681708930
transform 1 0 180 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1705
timestamp 1681708930
transform 1 0 180 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1776
timestamp 1681708930
transform 1 0 108 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1777
timestamp 1681708930
transform 1 0 164 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1778
timestamp 1681708930
transform 1 0 204 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1779
timestamp 1681708930
transform 1 0 260 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1780
timestamp 1681708930
transform 1 0 284 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1683
timestamp 1681708930
transform 1 0 164 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1648
timestamp 1681708930
transform 1 0 260 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_1839
timestamp 1681708930
transform 1 0 268 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_1649
timestamp 1681708930
transform 1 0 284 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_1781
timestamp 1681708930
transform 1 0 308 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1840
timestamp 1681708930
transform 1 0 300 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_1650
timestamp 1681708930
transform 1 0 308 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1593
timestamp 1681708930
transform 1 0 364 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1706
timestamp 1681708930
transform 1 0 364 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1782
timestamp 1681708930
transform 1 0 340 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1625
timestamp 1681708930
transform 1 0 364 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1566
timestamp 1681708930
transform 1 0 412 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1567
timestamp 1681708930
transform 1 0 460 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1568
timestamp 1681708930
transform 1 0 484 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1594
timestamp 1681708930
transform 1 0 428 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1707
timestamp 1681708930
transform 1 0 388 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1708
timestamp 1681708930
transform 1 0 476 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1709
timestamp 1681708930
transform 1 0 492 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1783
timestamp 1681708930
transform 1 0 380 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1784
timestamp 1681708930
transform 1 0 388 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1785
timestamp 1681708930
transform 1 0 428 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1841
timestamp 1681708930
transform 1 0 324 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1842
timestamp 1681708930
transform 1 0 332 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1843
timestamp 1681708930
transform 1 0 356 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1844
timestamp 1681708930
transform 1 0 364 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1857
timestamp 1681708930
transform 1 0 276 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_1684
timestamp 1681708930
transform 1 0 300 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_1858
timestamp 1681708930
transform 1 0 316 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_1685
timestamp 1681708930
transform 1 0 324 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_1859
timestamp 1681708930
transform 1 0 332 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_1626
timestamp 1681708930
transform 1 0 436 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1686
timestamp 1681708930
transform 1 0 412 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1541
timestamp 1681708930
transform 1 0 548 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1542
timestamp 1681708930
transform 1 0 596 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1569
timestamp 1681708930
transform 1 0 580 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1595
timestamp 1681708930
transform 1 0 540 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1710
timestamp 1681708930
transform 1 0 540 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1711
timestamp 1681708930
transform 1 0 548 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1712
timestamp 1681708930
transform 1 0 596 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1713
timestamp 1681708930
transform 1 0 604 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1786
timestamp 1681708930
transform 1 0 548 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1627
timestamp 1681708930
transform 1 0 564 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_1787
timestamp 1681708930
transform 1 0 604 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1651
timestamp 1681708930
transform 1 0 548 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1687
timestamp 1681708930
transform 1 0 604 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1596
timestamp 1681708930
transform 1 0 660 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1714
timestamp 1681708930
transform 1 0 652 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1715
timestamp 1681708930
transform 1 0 660 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_1628
timestamp 1681708930
transform 1 0 652 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1543
timestamp 1681708930
transform 1 0 716 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1544
timestamp 1681708930
transform 1 0 740 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1570
timestamp 1681708930
transform 1 0 716 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1597
timestamp 1681708930
transform 1 0 708 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1598
timestamp 1681708930
transform 1 0 740 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1545
timestamp 1681708930
transform 1 0 796 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_1716
timestamp 1681708930
transform 1 0 716 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1717
timestamp 1681708930
transform 1 0 740 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1718
timestamp 1681708930
transform 1 0 748 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1719
timestamp 1681708930
transform 1 0 756 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1788
timestamp 1681708930
transform 1 0 660 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1789
timestamp 1681708930
transform 1 0 684 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1790
timestamp 1681708930
transform 1 0 692 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1652
timestamp 1681708930
transform 1 0 692 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1688
timestamp 1681708930
transform 1 0 700 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1703
timestamp 1681708930
transform 1 0 684 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1715
timestamp 1681708930
transform 1 0 660 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_1791
timestamp 1681708930
transform 1 0 732 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1546
timestamp 1681708930
transform 1 0 828 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1571
timestamp 1681708930
transform 1 0 820 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1572
timestamp 1681708930
transform 1 0 852 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1599
timestamp 1681708930
transform 1 0 804 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1720
timestamp 1681708930
transform 1 0 804 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1721
timestamp 1681708930
transform 1 0 820 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1722
timestamp 1681708930
transform 1 0 836 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1723
timestamp 1681708930
transform 1 0 844 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_1629
timestamp 1681708930
transform 1 0 788 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1653
timestamp 1681708930
transform 1 0 748 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1630
timestamp 1681708930
transform 1 0 820 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_1792
timestamp 1681708930
transform 1 0 828 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1631
timestamp 1681708930
transform 1 0 844 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_1793
timestamp 1681708930
transform 1 0 852 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1654
timestamp 1681708930
transform 1 0 836 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1716
timestamp 1681708930
transform 1 0 804 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1547
timestamp 1681708930
transform 1 0 924 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1548
timestamp 1681708930
transform 1 0 956 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1573
timestamp 1681708930
transform 1 0 900 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1574
timestamp 1681708930
transform 1 0 972 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1600
timestamp 1681708930
transform 1 0 964 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1724
timestamp 1681708930
transform 1 0 876 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_1618
timestamp 1681708930
transform 1 0 900 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1601
timestamp 1681708930
transform 1 0 996 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1725
timestamp 1681708930
transform 1 0 964 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_1619
timestamp 1681708930
transform 1 0 972 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1575
timestamp 1681708930
transform 1 0 1020 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_1726
timestamp 1681708930
transform 1 0 980 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1727
timestamp 1681708930
transform 1 0 988 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1728
timestamp 1681708930
transform 1 0 1004 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1729
timestamp 1681708930
transform 1 0 1012 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1794
timestamp 1681708930
transform 1 0 860 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1795
timestamp 1681708930
transform 1 0 900 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1796
timestamp 1681708930
transform 1 0 956 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1797
timestamp 1681708930
transform 1 0 972 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1798
timestamp 1681708930
transform 1 0 980 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1799
timestamp 1681708930
transform 1 0 996 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1655
timestamp 1681708930
transform 1 0 860 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1656
timestamp 1681708930
transform 1 0 900 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1657
timestamp 1681708930
transform 1 0 916 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1658
timestamp 1681708930
transform 1 0 940 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1689
timestamp 1681708930
transform 1 0 852 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1717
timestamp 1681708930
transform 1 0 852 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1690
timestamp 1681708930
transform 1 0 956 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1718
timestamp 1681708930
transform 1 0 948 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1632
timestamp 1681708930
transform 1 0 1004 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1704
timestamp 1681708930
transform 1 0 980 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1633
timestamp 1681708930
transform 1 0 1028 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_1845
timestamp 1681708930
transform 1 0 1028 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_1549
timestamp 1681708930
transform 1 0 1108 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1550
timestamp 1681708930
transform 1 0 1124 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1551
timestamp 1681708930
transform 1 0 1148 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1552
timestamp 1681708930
transform 1 0 1180 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1553
timestamp 1681708930
transform 1 0 1212 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1576
timestamp 1681708930
transform 1 0 1060 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1577
timestamp 1681708930
transform 1 0 1100 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_1730
timestamp 1681708930
transform 1 0 1068 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1731
timestamp 1681708930
transform 1 0 1156 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1800
timestamp 1681708930
transform 1 0 1052 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1801
timestamp 1681708930
transform 1 0 1092 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1634
timestamp 1681708930
transform 1 0 1116 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1578
timestamp 1681708930
transform 1 0 1212 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1554
timestamp 1681708930
transform 1 0 1276 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1602
timestamp 1681708930
transform 1 0 1204 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1603
timestamp 1681708930
transform 1 0 1260 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1604
timestamp 1681708930
transform 1 0 1284 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1732
timestamp 1681708930
transform 1 0 1204 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1733
timestamp 1681708930
transform 1 0 1212 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1802
timestamp 1681708930
transform 1 0 1148 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1659
timestamp 1681708930
transform 1 0 1052 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1660
timestamp 1681708930
transform 1 0 1092 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1705
timestamp 1681708930
transform 1 0 1044 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1706
timestamp 1681708930
transform 1 0 1092 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1635
timestamp 1681708930
transform 1 0 1172 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_1803
timestamp 1681708930
transform 1 0 1180 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1804
timestamp 1681708930
transform 1 0 1204 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1691
timestamp 1681708930
transform 1 0 1164 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1719
timestamp 1681708930
transform 1 0 1068 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1720
timestamp 1681708930
transform 1 0 1148 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1636
timestamp 1681708930
transform 1 0 1268 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_1846
timestamp 1681708930
transform 1 0 1268 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_1555
timestamp 1681708930
transform 1 0 1308 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1605
timestamp 1681708930
transform 1 0 1308 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1606
timestamp 1681708930
transform 1 0 1340 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1734
timestamp 1681708930
transform 1 0 1292 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1735
timestamp 1681708930
transform 1 0 1308 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1736
timestamp 1681708930
transform 1 0 1316 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1805
timestamp 1681708930
transform 1 0 1300 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1661
timestamp 1681708930
transform 1 0 1292 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1620
timestamp 1681708930
transform 1 0 1324 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_1737
timestamp 1681708930
transform 1 0 1332 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1738
timestamp 1681708930
transform 1 0 1340 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_1621
timestamp 1681708930
transform 1 0 1356 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_1739
timestamp 1681708930
transform 1 0 1364 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1740
timestamp 1681708930
transform 1 0 1372 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1806
timestamp 1681708930
transform 1 0 1324 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1807
timestamp 1681708930
transform 1 0 1340 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1808
timestamp 1681708930
transform 1 0 1356 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1662
timestamp 1681708930
transform 1 0 1324 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1707
timestamp 1681708930
transform 1 0 1316 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1721
timestamp 1681708930
transform 1 0 1324 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_1809
timestamp 1681708930
transform 1 0 1380 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1556
timestamp 1681708930
transform 1 0 1404 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1607
timestamp 1681708930
transform 1 0 1404 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1608
timestamp 1681708930
transform 1 0 1436 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1741
timestamp 1681708930
transform 1 0 1404 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_1622
timestamp 1681708930
transform 1 0 1420 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_1742
timestamp 1681708930
transform 1 0 1428 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1743
timestamp 1681708930
transform 1 0 1436 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1810
timestamp 1681708930
transform 1 0 1396 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1811
timestamp 1681708930
transform 1 0 1404 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1812
timestamp 1681708930
transform 1 0 1420 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1813
timestamp 1681708930
transform 1 0 1436 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1663
timestamp 1681708930
transform 1 0 1396 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1664
timestamp 1681708930
transform 1 0 1436 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1692
timestamp 1681708930
transform 1 0 1428 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1708
timestamp 1681708930
transform 1 0 1404 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1557
timestamp 1681708930
transform 1 0 1524 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1609
timestamp 1681708930
transform 1 0 1508 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1701
timestamp 1681708930
transform 1 0 1516 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_1744
timestamp 1681708930
transform 1 0 1484 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1745
timestamp 1681708930
transform 1 0 1508 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1746
timestamp 1681708930
transform 1 0 1524 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_1637
timestamp 1681708930
transform 1 0 1460 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_1814
timestamp 1681708930
transform 1 0 1468 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1815
timestamp 1681708930
transform 1 0 1484 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1816
timestamp 1681708930
transform 1 0 1492 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1665
timestamp 1681708930
transform 1 0 1484 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_1817
timestamp 1681708930
transform 1 0 1524 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1666
timestamp 1681708930
transform 1 0 1524 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1709
timestamp 1681708930
transform 1 0 1500 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1638
timestamp 1681708930
transform 1 0 1540 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_1847
timestamp 1681708930
transform 1 0 1540 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_1693
timestamp 1681708930
transform 1 0 1540 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1610
timestamp 1681708930
transform 1 0 1564 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1747
timestamp 1681708930
transform 1 0 1564 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_1579
timestamp 1681708930
transform 1 0 1580 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_1848
timestamp 1681708930
transform 1 0 1572 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_1558
timestamp 1681708930
transform 1 0 1636 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_1748
timestamp 1681708930
transform 1 0 1612 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1849
timestamp 1681708930
transform 1 0 1596 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_1559
timestamp 1681708930
transform 1 0 1724 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1580
timestamp 1681708930
transform 1 0 1676 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_1749
timestamp 1681708930
transform 1 0 1668 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1750
timestamp 1681708930
transform 1 0 1716 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1751
timestamp 1681708930
transform 1 0 1724 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1818
timestamp 1681708930
transform 1 0 1628 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1860
timestamp 1681708930
transform 1 0 1604 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_1694
timestamp 1681708930
transform 1 0 1612 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1639
timestamp 1681708930
transform 1 0 1660 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1640
timestamp 1681708930
transform 1 0 1684 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1710
timestamp 1681708930
transform 1 0 1668 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1611
timestamp 1681708930
transform 1 0 1780 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1752
timestamp 1681708930
transform 1 0 1772 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1819
timestamp 1681708930
transform 1 0 1748 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1667
timestamp 1681708930
transform 1 0 1716 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1668
timestamp 1681708930
transform 1 0 1748 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1581
timestamp 1681708930
transform 1 0 1876 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_1753
timestamp 1681708930
transform 1 0 1828 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1754
timestamp 1681708930
transform 1 0 1836 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1820
timestamp 1681708930
transform 1 0 1804 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1641
timestamp 1681708930
transform 1 0 1828 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_1755
timestamp 1681708930
transform 1 0 1884 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1821
timestamp 1681708930
transform 1 0 1860 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1695
timestamp 1681708930
transform 1 0 1804 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1669
timestamp 1681708930
transform 1 0 1860 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1612
timestamp 1681708930
transform 1 0 1900 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1756
timestamp 1681708930
transform 1 0 1900 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_1560
timestamp 1681708930
transform 1 0 1932 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1582
timestamp 1681708930
transform 1 0 1916 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1583
timestamp 1681708930
transform 1 0 1972 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_1757
timestamp 1681708930
transform 1 0 1932 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1822
timestamp 1681708930
transform 1 0 1924 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1823
timestamp 1681708930
transform 1 0 1948 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1696
timestamp 1681708930
transform 1 0 1916 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1642
timestamp 1681708930
transform 1 0 1956 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1670
timestamp 1681708930
transform 1 0 1964 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1584
timestamp 1681708930
transform 1 0 2028 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_1758
timestamp 1681708930
transform 1 0 1996 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1759
timestamp 1681708930
transform 1 0 2004 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_1643
timestamp 1681708930
transform 1 0 1996 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_1824
timestamp 1681708930
transform 1 0 2004 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1697
timestamp 1681708930
transform 1 0 1996 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1671
timestamp 1681708930
transform 1 0 2052 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1722
timestamp 1681708930
transform 1 0 2020 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1561
timestamp 1681708930
transform 1 0 2076 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1613
timestamp 1681708930
transform 1 0 2068 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1672
timestamp 1681708930
transform 1 0 2068 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1562
timestamp 1681708930
transform 1 0 2100 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_1760
timestamp 1681708930
transform 1 0 2084 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1761
timestamp 1681708930
transform 1 0 2092 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_1698
timestamp 1681708930
transform 1 0 2084 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1723
timestamp 1681708930
transform 1 0 2076 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1585
timestamp 1681708930
transform 1 0 2140 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_1825
timestamp 1681708930
transform 1 0 2116 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1673
timestamp 1681708930
transform 1 0 2124 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1711
timestamp 1681708930
transform 1 0 2132 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_1762
timestamp 1681708930
transform 1 0 2148 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_1674
timestamp 1681708930
transform 1 0 2148 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1712
timestamp 1681708930
transform 1 0 2164 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_1763
timestamp 1681708930
transform 1 0 2180 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_1563
timestamp 1681708930
transform 1 0 2236 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1586
timestamp 1681708930
transform 1 0 2252 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1614
timestamp 1681708930
transform 1 0 2244 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1764
timestamp 1681708930
transform 1 0 2228 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1765
timestamp 1681708930
transform 1 0 2244 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1766
timestamp 1681708930
transform 1 0 2252 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1826
timestamp 1681708930
transform 1 0 2204 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1827
timestamp 1681708930
transform 1 0 2228 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1675
timestamp 1681708930
transform 1 0 2204 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1676
timestamp 1681708930
transform 1 0 2228 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1564
timestamp 1681708930
transform 1 0 2332 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_1767
timestamp 1681708930
transform 1 0 2300 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1768
timestamp 1681708930
transform 1 0 2308 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_1587
timestamp 1681708930
transform 1 0 2356 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_1769
timestamp 1681708930
transform 1 0 2356 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1828
timestamp 1681708930
transform 1 0 2324 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1829
timestamp 1681708930
transform 1 0 2332 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1830
timestamp 1681708930
transform 1 0 2356 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1699
timestamp 1681708930
transform 1 0 2356 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1615
timestamp 1681708930
transform 1 0 2380 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1850
timestamp 1681708930
transform 1 0 2380 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1770
timestamp 1681708930
transform 1 0 2388 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_1644
timestamp 1681708930
transform 1 0 2388 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1623
timestamp 1681708930
transform 1 0 2444 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_1831
timestamp 1681708930
transform 1 0 2412 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1645
timestamp 1681708930
transform 1 0 2428 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_1832
timestamp 1681708930
transform 1 0 2444 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1677
timestamp 1681708930
transform 1 0 2412 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1588
timestamp 1681708930
transform 1 0 2484 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1646
timestamp 1681708930
transform 1 0 2468 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_1833
timestamp 1681708930
transform 1 0 2476 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1851
timestamp 1681708930
transform 1 0 2420 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1852
timestamp 1681708930
transform 1 0 2428 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1861
timestamp 1681708930
transform 1 0 2404 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_1678
timestamp 1681708930
transform 1 0 2436 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_1853
timestamp 1681708930
transform 1 0 2444 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_1679
timestamp 1681708930
transform 1 0 2452 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_1854
timestamp 1681708930
transform 1 0 2460 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_1713
timestamp 1681708930
transform 1 0 2420 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_1855
timestamp 1681708930
transform 1 0 2484 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1862
timestamp 1681708930
transform 1 0 2452 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_1863
timestamp 1681708930
transform 1 0 2468 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_1864
timestamp 1681708930
transform 1 0 2476 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_1700
timestamp 1681708930
transform 1 0 2484 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1714
timestamp 1681708930
transform 1 0 2468 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1616
timestamp 1681708930
transform 1 0 2500 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1834
timestamp 1681708930
transform 1 0 2500 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1589
timestamp 1681708930
transform 1 0 2532 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1590
timestamp 1681708930
transform 1 0 2548 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_1702
timestamp 1681708930
transform 1 0 2516 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_1703
timestamp 1681708930
transform 1 0 2524 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_1624
timestamp 1681708930
transform 1 0 2524 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_1771
timestamp 1681708930
transform 1 0 2540 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1772
timestamp 1681708930
transform 1 0 2548 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1835
timestamp 1681708930
transform 1 0 2516 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1647
timestamp 1681708930
transform 1 0 2540 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1680
timestamp 1681708930
transform 1 0 2516 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1724
timestamp 1681708930
transform 1 0 2508 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_1836
timestamp 1681708930
transform 1 0 2564 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_1681
timestamp 1681708930
transform 1 0 2556 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1725
timestamp 1681708930
transform 1 0 2548 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1565
timestamp 1681708930
transform 1 0 2604 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1617
timestamp 1681708930
transform 1 0 2612 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_1773
timestamp 1681708930
transform 1 0 2604 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1774
timestamp 1681708930
transform 1 0 2612 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1837
timestamp 1681708930
transform 1 0 2588 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1838
timestamp 1681708930
transform 1 0 2596 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1856
timestamp 1681708930
transform 1 0 2572 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_1701
timestamp 1681708930
transform 1 0 2596 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_1775
timestamp 1681708930
transform 1 0 2732 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_1682
timestamp 1681708930
transform 1 0 2644 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1702
timestamp 1681708930
transform 1 0 2612 0 1 1505
box -3 -3 3 3
use top_mod_new_VIA0  top_mod_new_VIA0_22
timestamp 1681708930
transform 1 0 24 0 1 1470
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_36
timestamp 1681708930
transform 1 0 72 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_37
timestamp 1681708930
transform 1 0 168 0 -1 1570
box -8 -3 104 105
use NAND3X1  NAND3X1_61
timestamp 1681708930
transform -1 0 296 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_62
timestamp 1681708930
transform 1 0 296 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_63
timestamp 1681708930
transform 1 0 328 0 -1 1570
box -8 -3 40 105
use OAI21X1  OAI21X1_52
timestamp 1681708930
transform -1 0 392 0 -1 1570
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_38
timestamp 1681708930
transform -1 0 488 0 -1 1570
box -8 -3 104 105
use XNOR2X1  XNOR2X1_24
timestamp 1681708930
transform 1 0 488 0 -1 1570
box -8 -3 64 105
use XNOR2X1  XNOR2X1_26
timestamp 1681708930
transform 1 0 544 0 -1 1570
box -8 -3 64 105
use M3_M2  M3_M2_1726
timestamp 1681708930
transform 1 0 636 0 1 1475
box -3 -3 3 3
use XNOR2X1  XNOR2X1_27
timestamp 1681708930
transform 1 0 600 0 -1 1570
box -8 -3 64 105
use M3_M2  M3_M2_1727
timestamp 1681708930
transform 1 0 708 0 1 1475
box -3 -3 3 3
use XOR2X1  XOR2X1_65
timestamp 1681708930
transform 1 0 656 0 -1 1570
box -8 -3 64 105
use AOI22X1  AOI22X1_25
timestamp 1681708930
transform 1 0 712 0 -1 1570
box -8 -3 46 105
use XOR2X1  XOR2X1_66
timestamp 1681708930
transform 1 0 752 0 -1 1570
box -8 -3 64 105
use AOI22X1  AOI22X1_26
timestamp 1681708930
transform 1 0 808 0 -1 1570
box -8 -3 46 105
use INVX2  INVX2_109
timestamp 1681708930
transform 1 0 848 0 -1 1570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_41
timestamp 1681708930
transform 1 0 864 0 -1 1570
box -8 -3 104 105
use INVX2  INVX2_110
timestamp 1681708930
transform 1 0 960 0 -1 1570
box -9 -3 26 105
use M3_M2  M3_M2_1728
timestamp 1681708930
transform 1 0 1012 0 1 1475
box -3 -3 3 3
use AOI22X1  AOI22X1_27
timestamp 1681708930
transform 1 0 976 0 -1 1570
box -8 -3 46 105
use FILL  FILL_621
timestamp 1681708930
transform 1 0 1016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_622
timestamp 1681708930
transform 1 0 1024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_623
timestamp 1681708930
transform 1 0 1032 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_113
timestamp 1681708930
transform 1 0 1040 0 -1 1570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_42
timestamp 1681708930
transform 1 0 1056 0 -1 1570
box -8 -3 104 105
use M3_M2  M3_M2_1729
timestamp 1681708930
transform 1 0 1204 0 1 1475
box -3 -3 3 3
use XOR2X1  XOR2X1_74
timestamp 1681708930
transform -1 0 1208 0 -1 1570
box -8 -3 64 105
use XOR2X1  XOR2X1_75
timestamp 1681708930
transform -1 0 1264 0 -1 1570
box -8 -3 64 105
use OAI21X1  OAI21X1_53
timestamp 1681708930
transform -1 0 1296 0 -1 1570
box -8 -3 34 105
use NOR2X1  NOR2X1_43
timestamp 1681708930
transform 1 0 1296 0 -1 1570
box -8 -3 32 105
use INVX2  INVX2_114
timestamp 1681708930
transform -1 0 1336 0 -1 1570
box -9 -3 26 105
use AOI22X1  AOI22X1_29
timestamp 1681708930
transform 1 0 1336 0 -1 1570
box -8 -3 46 105
use FILL  FILL_644
timestamp 1681708930
transform 1 0 1376 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_115
timestamp 1681708930
transform 1 0 1384 0 -1 1570
box -9 -3 26 105
use AOI22X1  AOI22X1_30
timestamp 1681708930
transform 1 0 1400 0 -1 1570
box -8 -3 46 105
use FILL  FILL_645
timestamp 1681708930
transform 1 0 1440 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_31
timestamp 1681708930
transform -1 0 1488 0 -1 1570
box -8 -3 46 105
use OR2X1  OR2X1_10
timestamp 1681708930
transform -1 0 1520 0 -1 1570
box -8 -3 40 105
use NAND2X1  NAND2X1_49
timestamp 1681708930
transform 1 0 1520 0 -1 1570
box -8 -3 32 105
use INVX2  INVX2_116
timestamp 1681708930
transform -1 0 1560 0 -1 1570
box -9 -3 26 105
use FILL  FILL_646
timestamp 1681708930
transform 1 0 1560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_647
timestamp 1681708930
transform 1 0 1568 0 -1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_66
timestamp 1681708930
transform -1 0 1608 0 -1 1570
box -8 -3 40 105
use XNOR2X1  XNOR2X1_29
timestamp 1681708930
transform -1 0 1664 0 -1 1570
box -8 -3 64 105
use XOR2X1  XOR2X1_76
timestamp 1681708930
transform -1 0 1720 0 -1 1570
box -8 -3 64 105
use XOR2X1  XOR2X1_77
timestamp 1681708930
transform 1 0 1720 0 -1 1570
box -8 -3 64 105
use XOR2X1  XOR2X1_78
timestamp 1681708930
transform 1 0 1776 0 -1 1570
box -8 -3 64 105
use M3_M2  M3_M2_1730
timestamp 1681708930
transform 1 0 1884 0 1 1475
box -3 -3 3 3
use XOR2X1  XOR2X1_79
timestamp 1681708930
transform 1 0 1832 0 -1 1570
box -8 -3 64 105
use FILL  FILL_648
timestamp 1681708930
transform 1 0 1888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_649
timestamp 1681708930
transform 1 0 1896 0 -1 1570
box -8 -3 16 105
use FILL  FILL_651
timestamp 1681708930
transform 1 0 1904 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_117
timestamp 1681708930
transform 1 0 1912 0 -1 1570
box -9 -3 26 105
use XNOR2X1  XNOR2X1_30
timestamp 1681708930
transform -1 0 1984 0 -1 1570
box -8 -3 64 105
use FILL  FILL_659
timestamp 1681708930
transform 1 0 1984 0 -1 1570
box -8 -3 16 105
use FILL  FILL_660
timestamp 1681708930
transform 1 0 1992 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_1731
timestamp 1681708930
transform 1 0 2028 0 1 1475
box -3 -3 3 3
use XNOR2X1  XNOR2X1_31
timestamp 1681708930
transform -1 0 2056 0 -1 1570
box -8 -3 64 105
use FILL  FILL_661
timestamp 1681708930
transform 1 0 2056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_662
timestamp 1681708930
transform 1 0 2064 0 -1 1570
box -8 -3 16 105
use FILL  FILL_663
timestamp 1681708930
transform 1 0 2072 0 -1 1570
box -8 -3 16 105
use FILL  FILL_664
timestamp 1681708930
transform 1 0 2080 0 -1 1570
box -8 -3 16 105
use XOR2X1  XOR2X1_82
timestamp 1681708930
transform -1 0 2144 0 -1 1570
box -8 -3 64 105
use FILL  FILL_665
timestamp 1681708930
transform 1 0 2144 0 -1 1570
box -8 -3 16 105
use FILL  FILL_666
timestamp 1681708930
transform 1 0 2152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_667
timestamp 1681708930
transform 1 0 2160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_668
timestamp 1681708930
transform 1 0 2168 0 -1 1570
box -8 -3 16 105
use XOR2X1  XOR2X1_86
timestamp 1681708930
transform 1 0 2176 0 -1 1570
box -8 -3 64 105
use INVX2  INVX2_119
timestamp 1681708930
transform -1 0 2248 0 -1 1570
box -9 -3 26 105
use XOR2X1  XOR2X1_87
timestamp 1681708930
transform 1 0 2248 0 -1 1570
box -8 -3 64 105
use XOR2X1  XOR2X1_88
timestamp 1681708930
transform -1 0 2360 0 -1 1570
box -8 -3 64 105
use INVX2  INVX2_120
timestamp 1681708930
transform -1 0 2376 0 -1 1570
box -9 -3 26 105
use FILL  FILL_681
timestamp 1681708930
transform 1 0 2376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_682
timestamp 1681708930
transform 1 0 2384 0 -1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_70
timestamp 1681708930
transform -1 0 2424 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_71
timestamp 1681708930
transform -1 0 2456 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_72
timestamp 1681708930
transform -1 0 2488 0 -1 1570
box -8 -3 40 105
use FILL  FILL_683
timestamp 1681708930
transform 1 0 2488 0 -1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_45
timestamp 1681708930
transform -1 0 2520 0 -1 1570
box -8 -3 32 105
use AOI21X1  AOI21X1_29
timestamp 1681708930
transform -1 0 2552 0 -1 1570
box -7 -3 39 105
use FILL  FILL_684
timestamp 1681708930
transform 1 0 2552 0 -1 1570
box -8 -3 16 105
use FILL  FILL_685
timestamp 1681708930
transform 1 0 2560 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_54
timestamp 1681708930
transform -1 0 2600 0 -1 1570
box -8 -3 34 105
use FILL  FILL_686
timestamp 1681708930
transform 1 0 2600 0 -1 1570
box -8 -3 16 105
use XOR2X1  XOR2X1_89
timestamp 1681708930
transform -1 0 2664 0 -1 1570
box -8 -3 64 105
use top_mod_new_VIA0  top_mod_new_VIA0_23
timestamp 1681708930
transform 1 0 2712 0 1 1470
box -10 -3 10 3
use M3_M2  M3_M2_1755
timestamp 1681708930
transform 1 0 132 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_1865
timestamp 1681708930
transform 1 0 140 0 1 1435
box -2 -2 2 2
use M3_M2  M3_M2_1756
timestamp 1681708930
transform 1 0 156 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_1870
timestamp 1681708930
transform 1 0 132 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1871
timestamp 1681708930
transform 1 0 148 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1880
timestamp 1681708930
transform 1 0 132 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1797
timestamp 1681708930
transform 1 0 148 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_1872
timestamp 1681708930
transform 1 0 180 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1881
timestamp 1681708930
transform 1 0 156 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1882
timestamp 1681708930
transform 1 0 164 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1940
timestamp 1681708930
transform 1 0 156 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1798
timestamp 1681708930
transform 1 0 180 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1830
timestamp 1681708930
transform 1 0 156 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1831
timestamp 1681708930
transform 1 0 172 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_1941
timestamp 1681708930
transform 1 0 204 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2000
timestamp 1681708930
transform 1 0 220 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1942
timestamp 1681708930
transform 1 0 260 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1943
timestamp 1681708930
transform 1 0 268 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1944
timestamp 1681708930
transform 1 0 276 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1883
timestamp 1681708930
transform 1 0 292 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1945
timestamp 1681708930
transform 1 0 308 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1884
timestamp 1681708930
transform 1 0 340 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1866
timestamp 1681708930
transform 1 0 388 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_1873
timestamp 1681708930
transform 1 0 380 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1874
timestamp 1681708930
transform 1 0 404 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_1799
timestamp 1681708930
transform 1 0 380 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1800
timestamp 1681708930
transform 1 0 396 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_1946
timestamp 1681708930
transform 1 0 396 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1832
timestamp 1681708930
transform 1 0 396 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_1885
timestamp 1681708930
transform 1 0 428 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1947
timestamp 1681708930
transform 1 0 444 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1948
timestamp 1681708930
transform 1 0 452 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1833
timestamp 1681708930
transform 1 0 452 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_1886
timestamp 1681708930
transform 1 0 492 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1801
timestamp 1681708930
transform 1 0 532 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_1949
timestamp 1681708930
transform 1 0 500 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1850
timestamp 1681708930
transform 1 0 532 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1736
timestamp 1681708930
transform 1 0 556 0 1 1455
box -3 -3 3 3
use M2_M1  M2_M1_1887
timestamp 1681708930
transform 1 0 564 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1950
timestamp 1681708930
transform 1 0 556 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1802
timestamp 1681708930
transform 1 0 596 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_1951
timestamp 1681708930
transform 1 0 572 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1888
timestamp 1681708930
transform 1 0 628 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1952
timestamp 1681708930
transform 1 0 636 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1953
timestamp 1681708930
transform 1 0 644 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1771
timestamp 1681708930
transform 1 0 692 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_1889
timestamp 1681708930
transform 1 0 692 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1954
timestamp 1681708930
transform 1 0 700 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1955
timestamp 1681708930
transform 1 0 708 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2001
timestamp 1681708930
transform 1 0 700 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_1834
timestamp 1681708930
transform 1 0 708 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1803
timestamp 1681708930
transform 1 0 732 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1737
timestamp 1681708930
transform 1 0 756 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1757
timestamp 1681708930
transform 1 0 748 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1758
timestamp 1681708930
transform 1 0 764 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1759
timestamp 1681708930
transform 1 0 780 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1772
timestamp 1681708930
transform 1 0 756 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_1890
timestamp 1681708930
transform 1 0 748 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1891
timestamp 1681708930
transform 1 0 756 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1892
timestamp 1681708930
transform 1 0 772 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1804
timestamp 1681708930
transform 1 0 780 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_1893
timestamp 1681708930
transform 1 0 796 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1956
timestamp 1681708930
transform 1 0 756 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1957
timestamp 1681708930
transform 1 0 780 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1958
timestamp 1681708930
transform 1 0 788 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1835
timestamp 1681708930
transform 1 0 756 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1773
timestamp 1681708930
transform 1 0 828 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1760
timestamp 1681708930
transform 1 0 844 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1738
timestamp 1681708930
transform 1 0 868 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1761
timestamp 1681708930
transform 1 0 860 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_1894
timestamp 1681708930
transform 1 0 844 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1895
timestamp 1681708930
transform 1 0 852 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1959
timestamp 1681708930
transform 1 0 852 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1836
timestamp 1681708930
transform 1 0 852 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1744
timestamp 1681708930
transform 1 0 884 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1739
timestamp 1681708930
transform 1 0 916 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1745
timestamp 1681708930
transform 1 0 940 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1762
timestamp 1681708930
transform 1 0 924 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_1896
timestamp 1681708930
transform 1 0 900 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1805
timestamp 1681708930
transform 1 0 908 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_1897
timestamp 1681708930
transform 1 0 916 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1898
timestamp 1681708930
transform 1 0 924 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1960
timestamp 1681708930
transform 1 0 908 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1961
timestamp 1681708930
transform 1 0 916 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1763
timestamp 1681708930
transform 1 0 980 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1740
timestamp 1681708930
transform 1 0 1084 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1774
timestamp 1681708930
transform 1 0 1052 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_1899
timestamp 1681708930
transform 1 0 972 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1806
timestamp 1681708930
transform 1 0 996 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_1900
timestamp 1681708930
transform 1 0 1028 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1807
timestamp 1681708930
transform 1 0 1036 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_1901
timestamp 1681708930
transform 1 0 1052 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1962
timestamp 1681708930
transform 1 0 948 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1963
timestamp 1681708930
transform 1 0 1036 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1837
timestamp 1681708930
transform 1 0 932 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1838
timestamp 1681708930
transform 1 0 980 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1851
timestamp 1681708930
transform 1 0 1036 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1746
timestamp 1681708930
transform 1 0 1108 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1764
timestamp 1681708930
transform 1 0 1148 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1775
timestamp 1681708930
transform 1 0 1108 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1776
timestamp 1681708930
transform 1 0 1140 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1777
timestamp 1681708930
transform 1 0 1164 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1808
timestamp 1681708930
transform 1 0 1124 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_1902
timestamp 1681708930
transform 1 0 1140 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1903
timestamp 1681708930
transform 1 0 1148 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1964
timestamp 1681708930
transform 1 0 1084 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1965
timestamp 1681708930
transform 1 0 1092 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1839
timestamp 1681708930
transform 1 0 1084 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1809
timestamp 1681708930
transform 1 0 1172 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_1904
timestamp 1681708930
transform 1 0 1196 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1810
timestamp 1681708930
transform 1 0 1204 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_1905
timestamp 1681708930
transform 1 0 1220 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1966
timestamp 1681708930
transform 1 0 1140 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1967
timestamp 1681708930
transform 1 0 1148 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1840
timestamp 1681708930
transform 1 0 1140 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1747
timestamp 1681708930
transform 1 0 1244 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_1968
timestamp 1681708930
transform 1 0 1204 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1969
timestamp 1681708930
transform 1 0 1212 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1970
timestamp 1681708930
transform 1 0 1228 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1971
timestamp 1681708930
transform 1 0 1236 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1841
timestamp 1681708930
transform 1 0 1204 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1852
timestamp 1681708930
transform 1 0 1172 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1778
timestamp 1681708930
transform 1 0 1276 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_1906
timestamp 1681708930
transform 1 0 1260 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1907
timestamp 1681708930
transform 1 0 1268 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1842
timestamp 1681708930
transform 1 0 1260 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1748
timestamp 1681708930
transform 1 0 1308 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1765
timestamp 1681708930
transform 1 0 1300 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_1867
timestamp 1681708930
transform 1 0 1308 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_1875
timestamp 1681708930
transform 1 0 1292 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_1779
timestamp 1681708930
transform 1 0 1308 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_1908
timestamp 1681708930
transform 1 0 1300 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1821
timestamp 1681708930
transform 1 0 1300 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_1868
timestamp 1681708930
transform 1 0 1340 0 1 1435
box -2 -2 2 2
use M3_M2  M3_M2_1780
timestamp 1681708930
transform 1 0 1332 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_1876
timestamp 1681708930
transform 1 0 1348 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1909
timestamp 1681708930
transform 1 0 1332 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1843
timestamp 1681708930
transform 1 0 1316 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1811
timestamp 1681708930
transform 1 0 1348 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1741
timestamp 1681708930
transform 1 0 1364 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1749
timestamp 1681708930
transform 1 0 1372 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_1877
timestamp 1681708930
transform 1 0 1364 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_1781
timestamp 1681708930
transform 1 0 1404 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1750
timestamp 1681708930
transform 1 0 1452 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_1869
timestamp 1681708930
transform 1 0 1420 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_1878
timestamp 1681708930
transform 1 0 1412 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1910
timestamp 1681708930
transform 1 0 1404 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1822
timestamp 1681708930
transform 1 0 1388 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1766
timestamp 1681708930
transform 1 0 1428 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_1972
timestamp 1681708930
transform 1 0 1420 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1853
timestamp 1681708930
transform 1 0 1420 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_1911
timestamp 1681708930
transform 1 0 1436 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1912
timestamp 1681708930
transform 1 0 1452 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1823
timestamp 1681708930
transform 1 0 1436 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_1913
timestamp 1681708930
transform 1 0 1468 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1782
timestamp 1681708930
transform 1 0 1492 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1812
timestamp 1681708930
transform 1 0 1484 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_1973
timestamp 1681708930
transform 1 0 1444 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1974
timestamp 1681708930
transform 1 0 1460 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1824
timestamp 1681708930
transform 1 0 1468 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_1975
timestamp 1681708930
transform 1 0 1484 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1976
timestamp 1681708930
transform 1 0 1492 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1844
timestamp 1681708930
transform 1 0 1460 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_1914
timestamp 1681708930
transform 1 0 1500 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1845
timestamp 1681708930
transform 1 0 1500 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1783
timestamp 1681708930
transform 1 0 1532 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_1915
timestamp 1681708930
transform 1 0 1524 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1977
timestamp 1681708930
transform 1 0 1532 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1784
timestamp 1681708930
transform 1 0 1556 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_1916
timestamp 1681708930
transform 1 0 1564 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1767
timestamp 1681708930
transform 1 0 1580 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_1978
timestamp 1681708930
transform 1 0 1572 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1846
timestamp 1681708930
transform 1 0 1564 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1785
timestamp 1681708930
transform 1 0 1596 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1813
timestamp 1681708930
transform 1 0 1588 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_1917
timestamp 1681708930
transform 1 0 1612 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1979
timestamp 1681708930
transform 1 0 1596 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1980
timestamp 1681708930
transform 1 0 1604 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2002
timestamp 1681708930
transform 1 0 1580 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2003
timestamp 1681708930
transform 1 0 1612 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_1854
timestamp 1681708930
transform 1 0 1612 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1786
timestamp 1681708930
transform 1 0 1628 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_1918
timestamp 1681708930
transform 1 0 1628 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1751
timestamp 1681708930
transform 1 0 1644 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_1919
timestamp 1681708930
transform 1 0 1652 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1732
timestamp 1681708930
transform 1 0 1772 0 1 1465
box -3 -3 3 3
use M2_M1  M2_M1_1981
timestamp 1681708930
transform 1 0 1860 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1742
timestamp 1681708930
transform 1 0 1908 0 1 1455
box -3 -3 3 3
use M2_M1  M2_M1_1920
timestamp 1681708930
transform 1 0 1884 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1814
timestamp 1681708930
transform 1 0 1892 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_1921
timestamp 1681708930
transform 1 0 1900 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1922
timestamp 1681708930
transform 1 0 1916 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1825
timestamp 1681708930
transform 1 0 1884 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_1982
timestamp 1681708930
transform 1 0 1892 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1983
timestamp 1681708930
transform 1 0 1908 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1923
timestamp 1681708930
transform 1 0 1948 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1855
timestamp 1681708930
transform 1 0 1988 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_1924
timestamp 1681708930
transform 1 0 2004 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1733
timestamp 1681708930
transform 1 0 2052 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1752
timestamp 1681708930
transform 1 0 2052 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_1925
timestamp 1681708930
transform 1 0 2036 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1815
timestamp 1681708930
transform 1 0 2044 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_1926
timestamp 1681708930
transform 1 0 2052 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1984
timestamp 1681708930
transform 1 0 2044 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1985
timestamp 1681708930
transform 1 0 2052 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1856
timestamp 1681708930
transform 1 0 2036 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1753
timestamp 1681708930
transform 1 0 2164 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1768
timestamp 1681708930
transform 1 0 2132 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1787
timestamp 1681708930
transform 1 0 2068 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1788
timestamp 1681708930
transform 1 0 2108 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1769
timestamp 1681708930
transform 1 0 2196 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_1927
timestamp 1681708930
transform 1 0 2068 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1928
timestamp 1681708930
transform 1 0 2108 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1929
timestamp 1681708930
transform 1 0 2164 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1816
timestamp 1681708930
transform 1 0 2172 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1734
timestamp 1681708930
transform 1 0 2260 0 1 1465
box -3 -3 3 3
use M2_M1  M2_M1_1930
timestamp 1681708930
transform 1 0 2196 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1986
timestamp 1681708930
transform 1 0 2084 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1826
timestamp 1681708930
transform 1 0 2164 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_1987
timestamp 1681708930
transform 1 0 2172 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1857
timestamp 1681708930
transform 1 0 2148 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1817
timestamp 1681708930
transform 1 0 2220 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1743
timestamp 1681708930
transform 1 0 2276 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1754
timestamp 1681708930
transform 1 0 2284 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1789
timestamp 1681708930
transform 1 0 2276 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1790
timestamp 1681708930
transform 1 0 2308 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_1931
timestamp 1681708930
transform 1 0 2260 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1988
timestamp 1681708930
transform 1 0 2220 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1989
timestamp 1681708930
transform 1 0 2228 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1818
timestamp 1681708930
transform 1 0 2300 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_1932
timestamp 1681708930
transform 1 0 2308 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1990
timestamp 1681708930
transform 1 0 2276 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1991
timestamp 1681708930
transform 1 0 2284 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1847
timestamp 1681708930
transform 1 0 2276 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1858
timestamp 1681708930
transform 1 0 2244 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_1992
timestamp 1681708930
transform 1 0 2332 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1859
timestamp 1681708930
transform 1 0 2292 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1735
timestamp 1681708930
transform 1 0 2356 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1791
timestamp 1681708930
transform 1 0 2372 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1770
timestamp 1681708930
transform 1 0 2396 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_1993
timestamp 1681708930
transform 1 0 2388 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1933
timestamp 1681708930
transform 1 0 2404 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1934
timestamp 1681708930
transform 1 0 2444 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2004
timestamp 1681708930
transform 1 0 2436 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_1819
timestamp 1681708930
transform 1 0 2460 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1792
timestamp 1681708930
transform 1 0 2476 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_1879
timestamp 1681708930
transform 1 0 2484 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1935
timestamp 1681708930
transform 1 0 2476 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1994
timestamp 1681708930
transform 1 0 2460 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1995
timestamp 1681708930
transform 1 0 2468 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1848
timestamp 1681708930
transform 1 0 2452 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1820
timestamp 1681708930
transform 1 0 2484 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1793
timestamp 1681708930
transform 1 0 2516 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1827
timestamp 1681708930
transform 1 0 2508 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1794
timestamp 1681708930
transform 1 0 2532 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_1936
timestamp 1681708930
transform 1 0 2532 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1996
timestamp 1681708930
transform 1 0 2516 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1997
timestamp 1681708930
transform 1 0 2524 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1849
timestamp 1681708930
transform 1 0 2524 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_1937
timestamp 1681708930
transform 1 0 2548 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1828
timestamp 1681708930
transform 1 0 2540 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1795
timestamp 1681708930
transform 1 0 2564 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_1938
timestamp 1681708930
transform 1 0 2564 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_1829
timestamp 1681708930
transform 1 0 2556 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_1998
timestamp 1681708930
transform 1 0 2564 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1939
timestamp 1681708930
transform 1 0 2588 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1999
timestamp 1681708930
transform 1 0 2596 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_1796
timestamp 1681708930
transform 1 0 2628 0 1 1425
box -3 -3 3 3
use top_mod_new_VIA0  top_mod_new_VIA0_24
timestamp 1681708930
transform 1 0 48 0 1 1370
box -10 -3 10 3
use FILL  FILL_687
timestamp 1681708930
transform 1 0 72 0 1 1370
box -8 -3 16 105
use FILL  FILL_689
timestamp 1681708930
transform 1 0 80 0 1 1370
box -8 -3 16 105
use FILL  FILL_691
timestamp 1681708930
transform 1 0 88 0 1 1370
box -8 -3 16 105
use FILL  FILL_693
timestamp 1681708930
transform 1 0 96 0 1 1370
box -8 -3 16 105
use FILL  FILL_695
timestamp 1681708930
transform 1 0 104 0 1 1370
box -8 -3 16 105
use FILL  FILL_696
timestamp 1681708930
transform 1 0 112 0 1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_73
timestamp 1681708930
transform 1 0 120 0 1 1370
box -8 -3 40 105
use OAI21X1  OAI21X1_55
timestamp 1681708930
transform 1 0 152 0 1 1370
box -8 -3 34 105
use FILL  FILL_697
timestamp 1681708930
transform 1 0 184 0 1 1370
box -8 -3 16 105
use FILL  FILL_698
timestamp 1681708930
transform 1 0 192 0 1 1370
box -8 -3 16 105
use FILL  FILL_699
timestamp 1681708930
transform 1 0 200 0 1 1370
box -8 -3 16 105
use FILL  FILL_700
timestamp 1681708930
transform 1 0 208 0 1 1370
box -8 -3 16 105
use FILL  FILL_701
timestamp 1681708930
transform 1 0 216 0 1 1370
box -8 -3 16 105
use FILL  FILL_702
timestamp 1681708930
transform 1 0 224 0 1 1370
box -8 -3 16 105
use FILL  FILL_703
timestamp 1681708930
transform 1 0 232 0 1 1370
box -8 -3 16 105
use FILL  FILL_704
timestamp 1681708930
transform 1 0 240 0 1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_46
timestamp 1681708930
transform 1 0 248 0 1 1370
box -8 -3 32 105
use INVX2  INVX2_121
timestamp 1681708930
transform 1 0 272 0 1 1370
box -9 -3 26 105
use FILL  FILL_705
timestamp 1681708930
transform 1 0 288 0 1 1370
box -8 -3 16 105
use FILL  FILL_706
timestamp 1681708930
transform 1 0 296 0 1 1370
box -8 -3 16 105
use FILL  FILL_707
timestamp 1681708930
transform 1 0 304 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_122
timestamp 1681708930
transform 1 0 312 0 1 1370
box -9 -3 26 105
use FILL  FILL_708
timestamp 1681708930
transform 1 0 328 0 1 1370
box -8 -3 16 105
use FILL  FILL_709
timestamp 1681708930
transform 1 0 336 0 1 1370
box -8 -3 16 105
use FILL  FILL_710
timestamp 1681708930
transform 1 0 344 0 1 1370
box -8 -3 16 105
use FILL  FILL_715
timestamp 1681708930
transform 1 0 352 0 1 1370
box -8 -3 16 105
use FILL  FILL_717
timestamp 1681708930
transform 1 0 360 0 1 1370
box -8 -3 16 105
use FILL  FILL_719
timestamp 1681708930
transform 1 0 368 0 1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_75
timestamp 1681708930
transform -1 0 408 0 1 1370
box -8 -3 40 105
use FILL  FILL_720
timestamp 1681708930
transform 1 0 408 0 1 1370
box -8 -3 16 105
use FILL  FILL_721
timestamp 1681708930
transform 1 0 416 0 1 1370
box -8 -3 16 105
use BUFX2  BUFX2_3
timestamp 1681708930
transform 1 0 424 0 1 1370
box -5 -3 28 105
use FILL  FILL_722
timestamp 1681708930
transform 1 0 448 0 1 1370
box -8 -3 16 105
use FILL  FILL_723
timestamp 1681708930
transform 1 0 456 0 1 1370
box -8 -3 16 105
use FILL  FILL_724
timestamp 1681708930
transform 1 0 464 0 1 1370
box -8 -3 16 105
use FILL  FILL_725
timestamp 1681708930
transform 1 0 472 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_125
timestamp 1681708930
transform 1 0 480 0 1 1370
box -9 -3 26 105
use XOR2X1  XOR2X1_90
timestamp 1681708930
transform 1 0 496 0 1 1370
box -8 -3 64 105
use FILL  FILL_726
timestamp 1681708930
transform 1 0 552 0 1 1370
box -8 -3 16 105
use FILL  FILL_734
timestamp 1681708930
transform 1 0 560 0 1 1370
box -8 -3 16 105
use XOR2X1  XOR2X1_92
timestamp 1681708930
transform 1 0 568 0 1 1370
box -8 -3 64 105
use FILL  FILL_736
timestamp 1681708930
transform 1 0 624 0 1 1370
box -8 -3 16 105
use FILL  FILL_741
timestamp 1681708930
transform 1 0 632 0 1 1370
box -8 -3 16 105
use XOR2X1  XOR2X1_93
timestamp 1681708930
transform 1 0 640 0 1 1370
box -8 -3 64 105
use OR2X1  OR2X1_11
timestamp 1681708930
transform 1 0 696 0 1 1370
box -8 -3 40 105
use FILL  FILL_743
timestamp 1681708930
transform 1 0 728 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_127
timestamp 1681708930
transform 1 0 736 0 1 1370
box -9 -3 26 105
use AOI22X1  AOI22X1_32
timestamp 1681708930
transform 1 0 752 0 1 1370
box -8 -3 46 105
use FILL  FILL_756
timestamp 1681708930
transform 1 0 792 0 1 1370
box -8 -3 16 105
use FILL  FILL_757
timestamp 1681708930
transform 1 0 800 0 1 1370
box -8 -3 16 105
use FILL  FILL_758
timestamp 1681708930
transform 1 0 808 0 1 1370
box -8 -3 16 105
use FILL  FILL_759
timestamp 1681708930
transform 1 0 816 0 1 1370
box -8 -3 16 105
use FILL  FILL_760
timestamp 1681708930
transform 1 0 824 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_128
timestamp 1681708930
transform 1 0 832 0 1 1370
box -9 -3 26 105
use FILL  FILL_761
timestamp 1681708930
transform 1 0 848 0 1 1370
box -8 -3 16 105
use FILL  FILL_762
timestamp 1681708930
transform 1 0 856 0 1 1370
box -8 -3 16 105
use FILL  FILL_763
timestamp 1681708930
transform 1 0 864 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_1860
timestamp 1681708930
transform 1 0 892 0 1 1375
box -3 -3 3 3
use FILL  FILL_764
timestamp 1681708930
transform 1 0 872 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_33
timestamp 1681708930
transform 1 0 880 0 1 1370
box -8 -3 46 105
use INVX2  INVX2_129
timestamp 1681708930
transform 1 0 920 0 1 1370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_45
timestamp 1681708930
transform 1 0 936 0 1 1370
box -8 -3 104 105
use XOR2X1  XOR2X1_94
timestamp 1681708930
transform -1 0 1088 0 1 1370
box -8 -3 64 105
use M3_M2  M3_M2_1861
timestamp 1681708930
transform 1 0 1100 0 1 1375
box -3 -3 3 3
use XOR2X1  XOR2X1_95
timestamp 1681708930
transform 1 0 1088 0 1 1370
box -8 -3 64 105
use M3_M2  M3_M2_1862
timestamp 1681708930
transform 1 0 1156 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1863
timestamp 1681708930
transform 1 0 1172 0 1 1375
box -3 -3 3 3
use XOR2X1  XOR2X1_96
timestamp 1681708930
transform -1 0 1200 0 1 1370
box -8 -3 64 105
use M3_M2  M3_M2_1864
timestamp 1681708930
transform 1 0 1252 0 1 1375
box -3 -3 3 3
use AOI22X1  AOI22X1_34
timestamp 1681708930
transform 1 0 1200 0 1 1370
box -8 -3 46 105
use FILL  FILL_765
timestamp 1681708930
transform 1 0 1240 0 1 1370
box -8 -3 16 105
use FILL  FILL_766
timestamp 1681708930
transform 1 0 1248 0 1 1370
box -8 -3 16 105
use FILL  FILL_767
timestamp 1681708930
transform 1 0 1256 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_130
timestamp 1681708930
transform 1 0 1264 0 1 1370
box -9 -3 26 105
use FILL  FILL_768
timestamp 1681708930
transform 1 0 1280 0 1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_79
timestamp 1681708930
transform 1 0 1288 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_80
timestamp 1681708930
transform 1 0 1320 0 1 1370
box -8 -3 40 105
use FILL  FILL_769
timestamp 1681708930
transform 1 0 1352 0 1 1370
box -8 -3 16 105
use FILL  FILL_770
timestamp 1681708930
transform 1 0 1360 0 1 1370
box -8 -3 16 105
use FILL  FILL_771
timestamp 1681708930
transform 1 0 1368 0 1 1370
box -8 -3 16 105
use FILL  FILL_772
timestamp 1681708930
transform 1 0 1376 0 1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_81
timestamp 1681708930
transform -1 0 1416 0 1 1370
box -8 -3 40 105
use FILL  FILL_773
timestamp 1681708930
transform 1 0 1416 0 1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_21
timestamp 1681708930
transform 1 0 1424 0 1 1370
box -8 -3 46 105
use FILL  FILL_774
timestamp 1681708930
transform 1 0 1464 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_1865
timestamp 1681708930
transform 1 0 1484 0 1 1375
box -3 -3 3 3
use INVX2  INVX2_131
timestamp 1681708930
transform -1 0 1488 0 1 1370
box -9 -3 26 105
use M3_M2  M3_M2_1866
timestamp 1681708930
transform 1 0 1500 0 1 1375
box -3 -3 3 3
use FILL  FILL_775
timestamp 1681708930
transform 1 0 1488 0 1 1370
box -8 -3 16 105
use FILL  FILL_776
timestamp 1681708930
transform 1 0 1496 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_1867
timestamp 1681708930
transform 1 0 1516 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1868
timestamp 1681708930
transform 1 0 1540 0 1 1375
box -3 -3 3 3
use AOI22X1  AOI22X1_35
timestamp 1681708930
transform 1 0 1504 0 1 1370
box -8 -3 46 105
use INVX2  INVX2_132
timestamp 1681708930
transform -1 0 1560 0 1 1370
box -9 -3 26 105
use FILL  FILL_777
timestamp 1681708930
transform 1 0 1560 0 1 1370
box -8 -3 16 105
use FILL  FILL_778
timestamp 1681708930
transform 1 0 1568 0 1 1370
box -8 -3 16 105
use AOI21X1  AOI21X1_31
timestamp 1681708930
transform -1 0 1608 0 1 1370
box -7 -3 39 105
use NOR2X1  NOR2X1_48
timestamp 1681708930
transform 1 0 1608 0 1 1370
box -8 -3 32 105
use FILL  FILL_779
timestamp 1681708930
transform 1 0 1632 0 1 1370
box -8 -3 16 105
use FILL  FILL_780
timestamp 1681708930
transform 1 0 1640 0 1 1370
box -8 -3 16 105
use FILL  FILL_781
timestamp 1681708930
transform 1 0 1648 0 1 1370
box -8 -3 16 105
use FILL  FILL_782
timestamp 1681708930
transform 1 0 1656 0 1 1370
box -8 -3 16 105
use FILL  FILL_783
timestamp 1681708930
transform 1 0 1664 0 1 1370
box -8 -3 16 105
use FILL  FILL_784
timestamp 1681708930
transform 1 0 1672 0 1 1370
box -8 -3 16 105
use FILL  FILL_785
timestamp 1681708930
transform 1 0 1680 0 1 1370
box -8 -3 16 105
use FILL  FILL_786
timestamp 1681708930
transform 1 0 1688 0 1 1370
box -8 -3 16 105
use FILL  FILL_787
timestamp 1681708930
transform 1 0 1696 0 1 1370
box -8 -3 16 105
use FILL  FILL_788
timestamp 1681708930
transform 1 0 1704 0 1 1370
box -8 -3 16 105
use FILL  FILL_789
timestamp 1681708930
transform 1 0 1712 0 1 1370
box -8 -3 16 105
use FILL  FILL_790
timestamp 1681708930
transform 1 0 1720 0 1 1370
box -8 -3 16 105
use FILL  FILL_791
timestamp 1681708930
transform 1 0 1728 0 1 1370
box -8 -3 16 105
use FILL  FILL_792
timestamp 1681708930
transform 1 0 1736 0 1 1370
box -8 -3 16 105
use FILL  FILL_793
timestamp 1681708930
transform 1 0 1744 0 1 1370
box -8 -3 16 105
use FILL  FILL_794
timestamp 1681708930
transform 1 0 1752 0 1 1370
box -8 -3 16 105
use FILL  FILL_795
timestamp 1681708930
transform 1 0 1760 0 1 1370
box -8 -3 16 105
use FILL  FILL_796
timestamp 1681708930
transform 1 0 1768 0 1 1370
box -8 -3 16 105
use FILL  FILL_797
timestamp 1681708930
transform 1 0 1776 0 1 1370
box -8 -3 16 105
use FILL  FILL_798
timestamp 1681708930
transform 1 0 1784 0 1 1370
box -8 -3 16 105
use FILL  FILL_799
timestamp 1681708930
transform 1 0 1792 0 1 1370
box -8 -3 16 105
use FILL  FILL_800
timestamp 1681708930
transform 1 0 1800 0 1 1370
box -8 -3 16 105
use FILL  FILL_801
timestamp 1681708930
transform 1 0 1808 0 1 1370
box -8 -3 16 105
use FILL  FILL_802
timestamp 1681708930
transform 1 0 1816 0 1 1370
box -8 -3 16 105
use FILL  FILL_803
timestamp 1681708930
transform 1 0 1824 0 1 1370
box -8 -3 16 105
use FILL  FILL_804
timestamp 1681708930
transform 1 0 1832 0 1 1370
box -8 -3 16 105
use FILL  FILL_828
timestamp 1681708930
transform 1 0 1840 0 1 1370
box -8 -3 16 105
use FILL  FILL_830
timestamp 1681708930
transform 1 0 1848 0 1 1370
box -8 -3 16 105
use FILL  FILL_832
timestamp 1681708930
transform 1 0 1856 0 1 1370
box -8 -3 16 105
use FILL  FILL_833
timestamp 1681708930
transform 1 0 1864 0 1 1370
box -8 -3 16 105
use FILL  FILL_834
timestamp 1681708930
transform 1 0 1872 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_43
timestamp 1681708930
transform -1 0 1920 0 1 1370
box -8 -3 46 105
use FILL  FILL_835
timestamp 1681708930
transform 1 0 1920 0 1 1370
box -8 -3 16 105
use FILL  FILL_836
timestamp 1681708930
transform 1 0 1928 0 1 1370
box -8 -3 16 105
use FILL  FILL_837
timestamp 1681708930
transform 1 0 1936 0 1 1370
box -8 -3 16 105
use FILL  FILL_838
timestamp 1681708930
transform 1 0 1944 0 1 1370
box -8 -3 16 105
use FILL  FILL_839
timestamp 1681708930
transform 1 0 1952 0 1 1370
box -8 -3 16 105
use FILL  FILL_840
timestamp 1681708930
transform 1 0 1960 0 1 1370
box -8 -3 16 105
use FILL  FILL_841
timestamp 1681708930
transform 1 0 1968 0 1 1370
box -8 -3 16 105
use FILL  FILL_842
timestamp 1681708930
transform 1 0 1976 0 1 1370
box -8 -3 16 105
use FILL  FILL_843
timestamp 1681708930
transform 1 0 1984 0 1 1370
box -8 -3 16 105
use FILL  FILL_844
timestamp 1681708930
transform 1 0 1992 0 1 1370
box -8 -3 16 105
use FILL  FILL_845
timestamp 1681708930
transform 1 0 2000 0 1 1370
box -8 -3 16 105
use FILL  FILL_846
timestamp 1681708930
transform 1 0 2008 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_1869
timestamp 1681708930
transform 1 0 2028 0 1 1375
box -3 -3 3 3
use AOI22X1  AOI22X1_44
timestamp 1681708930
transform 1 0 2016 0 1 1370
box -8 -3 46 105
use INVX2  INVX2_139
timestamp 1681708930
transform 1 0 2056 0 1 1370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_50
timestamp 1681708930
transform 1 0 2072 0 1 1370
box -8 -3 104 105
use XOR2X1  XOR2X1_98
timestamp 1681708930
transform -1 0 2224 0 1 1370
box -8 -3 64 105
use M3_M2  M3_M2_1870
timestamp 1681708930
transform 1 0 2244 0 1 1375
box -3 -3 3 3
use XOR2X1  XOR2X1_99
timestamp 1681708930
transform 1 0 2224 0 1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_100
timestamp 1681708930
transform -1 0 2336 0 1 1370
box -8 -3 64 105
use FILL  FILL_847
timestamp 1681708930
transform 1 0 2336 0 1 1370
box -8 -3 16 105
use FILL  FILL_848
timestamp 1681708930
transform 1 0 2344 0 1 1370
box -8 -3 16 105
use FILL  FILL_849
timestamp 1681708930
transform 1 0 2352 0 1 1370
box -8 -3 16 105
use FILL  FILL_850
timestamp 1681708930
transform 1 0 2360 0 1 1370
box -8 -3 16 105
use FILL  FILL_851
timestamp 1681708930
transform 1 0 2368 0 1 1370
box -8 -3 16 105
use FILL  FILL_852
timestamp 1681708930
transform 1 0 2376 0 1 1370
box -8 -3 16 105
use FILL  FILL_853
timestamp 1681708930
transform 1 0 2384 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_140
timestamp 1681708930
transform 1 0 2392 0 1 1370
box -9 -3 26 105
use FILL  FILL_854
timestamp 1681708930
transform 1 0 2408 0 1 1370
box -8 -3 16 105
use FILL  FILL_855
timestamp 1681708930
transform 1 0 2416 0 1 1370
box -8 -3 16 105
use FILL  FILL_856
timestamp 1681708930
transform 1 0 2424 0 1 1370
box -8 -3 16 105
use FILL  FILL_857
timestamp 1681708930
transform 1 0 2432 0 1 1370
box -8 -3 16 105
use AOI21X1  AOI21X1_32
timestamp 1681708930
transform -1 0 2472 0 1 1370
box -7 -3 39 105
use FILL  FILL_858
timestamp 1681708930
transform 1 0 2472 0 1 1370
box -8 -3 16 105
use FILL  FILL_859
timestamp 1681708930
transform 1 0 2480 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_57
timestamp 1681708930
transform -1 0 2520 0 1 1370
box -8 -3 34 105
use FILL  FILL_860
timestamp 1681708930
transform 1 0 2520 0 1 1370
box -8 -3 16 105
use FILL  FILL_861
timestamp 1681708930
transform 1 0 2528 0 1 1370
box -8 -3 16 105
use FILL  FILL_862
timestamp 1681708930
transform 1 0 2536 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_141
timestamp 1681708930
transform 1 0 2544 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_142
timestamp 1681708930
transform 1 0 2560 0 1 1370
box -9 -3 26 105
use NAND2X1  NAND2X1_52
timestamp 1681708930
transform -1 0 2600 0 1 1370
box -8 -3 32 105
use FILL  FILL_863
timestamp 1681708930
transform 1 0 2600 0 1 1370
box -8 -3 16 105
use FILL  FILL_864
timestamp 1681708930
transform 1 0 2608 0 1 1370
box -8 -3 16 105
use FILL  FILL_865
timestamp 1681708930
transform 1 0 2616 0 1 1370
box -8 -3 16 105
use FILL  FILL_866
timestamp 1681708930
transform 1 0 2624 0 1 1370
box -8 -3 16 105
use FILL  FILL_867
timestamp 1681708930
transform 1 0 2632 0 1 1370
box -8 -3 16 105
use FILL  FILL_871
timestamp 1681708930
transform 1 0 2640 0 1 1370
box -8 -3 16 105
use FILL  FILL_873
timestamp 1681708930
transform 1 0 2648 0 1 1370
box -8 -3 16 105
use FILL  FILL_875
timestamp 1681708930
transform 1 0 2656 0 1 1370
box -8 -3 16 105
use top_mod_new_VIA0  top_mod_new_VIA0_25
timestamp 1681708930
transform 1 0 2688 0 1 1370
box -10 -3 10 3
use M2_M1  M2_M1_2075
timestamp 1681708930
transform 1 0 100 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2005
timestamp 1681708930
transform 1 0 108 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2012
timestamp 1681708930
transform 1 0 132 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_1948
timestamp 1681708930
transform 1 0 132 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_2076
timestamp 1681708930
transform 1 0 140 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2077
timestamp 1681708930
transform 1 0 148 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1907
timestamp 1681708930
transform 1 0 156 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_2013
timestamp 1681708930
transform 1 0 156 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2078
timestamp 1681708930
transform 1 0 156 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1908
timestamp 1681708930
transform 1 0 220 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_2014
timestamp 1681708930
transform 1 0 172 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2015
timestamp 1681708930
transform 1 0 188 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_1933
timestamp 1681708930
transform 1 0 268 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_2079
timestamp 1681708930
transform 1 0 212 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2080
timestamp 1681708930
transform 1 0 268 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1968
timestamp 1681708930
transform 1 0 220 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1997
timestamp 1681708930
transform 1 0 180 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1998
timestamp 1681708930
transform 1 0 212 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2025
timestamp 1681708930
transform 1 0 172 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1949
timestamp 1681708930
transform 1 0 276 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_2006
timestamp 1681708930
transform 1 0 292 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_1909
timestamp 1681708930
transform 1 0 300 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1934
timestamp 1681708930
transform 1 0 292 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_2016
timestamp 1681708930
transform 1 0 300 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2017
timestamp 1681708930
transform 1 0 308 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_2017
timestamp 1681708930
transform 1 0 284 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2026
timestamp 1681708930
transform 1 0 284 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1935
timestamp 1681708930
transform 1 0 316 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_2018
timestamp 1681708930
transform 1 0 324 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_1950
timestamp 1681708930
transform 1 0 316 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_2144
timestamp 1681708930
transform 1 0 316 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2159
timestamp 1681708930
transform 1 0 316 0 1 1305
box -2 -2 2 2
use M3_M2  M3_M2_2018
timestamp 1681708930
transform 1 0 300 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1910
timestamp 1681708930
transform 1 0 348 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_2019
timestamp 1681708930
transform 1 0 348 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2081
timestamp 1681708930
transform 1 0 356 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2020
timestamp 1681708930
transform 1 0 372 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_1951
timestamp 1681708930
transform 1 0 364 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_2145
timestamp 1681708930
transform 1 0 364 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_1952
timestamp 1681708930
transform 1 0 396 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1871
timestamp 1681708930
transform 1 0 412 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1884
timestamp 1681708930
transform 1 0 428 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_2021
timestamp 1681708930
transform 1 0 412 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_1885
timestamp 1681708930
transform 1 0 484 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_2022
timestamp 1681708930
transform 1 0 460 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2082
timestamp 1681708930
transform 1 0 428 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2083
timestamp 1681708930
transform 1 0 476 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2146
timestamp 1681708930
transform 1 0 468 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_1969
timestamp 1681708930
transform 1 0 476 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1999
timestamp 1681708930
transform 1 0 444 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2000
timestamp 1681708930
transform 1 0 468 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_2160
timestamp 1681708930
transform 1 0 476 0 1 1305
box -2 -2 2 2
use M3_M2  M3_M2_1936
timestamp 1681708930
transform 1 0 524 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_2084
timestamp 1681708930
transform 1 0 524 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2147
timestamp 1681708930
transform 1 0 500 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2148
timestamp 1681708930
transform 1 0 508 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2149
timestamp 1681708930
transform 1 0 524 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2001
timestamp 1681708930
transform 1 0 500 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_2161
timestamp 1681708930
transform 1 0 516 0 1 1305
box -2 -2 2 2
use M3_M2  M3_M2_2002
timestamp 1681708930
transform 1 0 524 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_2150
timestamp 1681708930
transform 1 0 572 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2003
timestamp 1681708930
transform 1 0 572 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1937
timestamp 1681708930
transform 1 0 604 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_2085
timestamp 1681708930
transform 1 0 604 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2151
timestamp 1681708930
transform 1 0 612 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2162
timestamp 1681708930
transform 1 0 596 0 1 1305
box -2 -2 2 2
use M3_M2  M3_M2_1872
timestamp 1681708930
transform 1 0 644 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1911
timestamp 1681708930
transform 1 0 700 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_2086
timestamp 1681708930
transform 1 0 692 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2023
timestamp 1681708930
transform 1 0 708 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2024
timestamp 1681708930
transform 1 0 764 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_1953
timestamp 1681708930
transform 1 0 740 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1873
timestamp 1681708930
transform 1 0 780 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_2087
timestamp 1681708930
transform 1 0 756 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2088
timestamp 1681708930
transform 1 0 772 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1886
timestamp 1681708930
transform 1 0 788 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1874
timestamp 1681708930
transform 1 0 820 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1875
timestamp 1681708930
transform 1 0 868 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1876
timestamp 1681708930
transform 1 0 884 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1912
timestamp 1681708930
transform 1 0 876 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_2025
timestamp 1681708930
transform 1 0 876 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2089
timestamp 1681708930
transform 1 0 796 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2090
timestamp 1681708930
transform 1 0 844 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2004
timestamp 1681708930
transform 1 0 796 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2019
timestamp 1681708930
transform 1 0 804 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2027
timestamp 1681708930
transform 1 0 804 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1913
timestamp 1681708930
transform 1 0 900 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1914
timestamp 1681708930
transform 1 0 948 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_2026
timestamp 1681708930
transform 1 0 900 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_1887
timestamp 1681708930
transform 1 0 988 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_2091
timestamp 1681708930
transform 1 0 924 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2092
timestamp 1681708930
transform 1 0 980 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1915
timestamp 1681708930
transform 1 0 996 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_2027
timestamp 1681708930
transform 1 0 996 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2093
timestamp 1681708930
transform 1 0 1004 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1970
timestamp 1681708930
transform 1 0 996 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1877
timestamp 1681708930
transform 1 0 1044 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1888
timestamp 1681708930
transform 1 0 1028 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_2028
timestamp 1681708930
transform 1 0 1028 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_1938
timestamp 1681708930
transform 1 0 1036 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_2094
timestamp 1681708930
transform 1 0 1020 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2095
timestamp 1681708930
transform 1 0 1036 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1971
timestamp 1681708930
transform 1 0 1036 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_2096
timestamp 1681708930
transform 1 0 1060 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1889
timestamp 1681708930
transform 1 0 1076 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1916
timestamp 1681708930
transform 1 0 1068 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_2029
timestamp 1681708930
transform 1 0 1068 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2030
timestamp 1681708930
transform 1 0 1076 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2097
timestamp 1681708930
transform 1 0 1084 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2020
timestamp 1681708930
transform 1 0 1084 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1890
timestamp 1681708930
transform 1 0 1132 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1917
timestamp 1681708930
transform 1 0 1124 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_2031
timestamp 1681708930
transform 1 0 1124 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2032
timestamp 1681708930
transform 1 0 1132 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2098
timestamp 1681708930
transform 1 0 1116 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2099
timestamp 1681708930
transform 1 0 1148 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2100
timestamp 1681708930
transform 1 0 1156 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1878
timestamp 1681708930
transform 1 0 1172 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1891
timestamp 1681708930
transform 1 0 1180 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1918
timestamp 1681708930
transform 1 0 1196 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_2033
timestamp 1681708930
transform 1 0 1180 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2034
timestamp 1681708930
transform 1 0 1196 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2101
timestamp 1681708930
transform 1 0 1188 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1892
timestamp 1681708930
transform 1 0 1212 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_2102
timestamp 1681708930
transform 1 0 1212 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1919
timestamp 1681708930
transform 1 0 1220 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1939
timestamp 1681708930
transform 1 0 1220 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1972
timestamp 1681708930
transform 1 0 1212 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1879
timestamp 1681708930
transform 1 0 1244 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1880
timestamp 1681708930
transform 1 0 1324 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_2035
timestamp 1681708930
transform 1 0 1236 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2036
timestamp 1681708930
transform 1 0 1324 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2103
timestamp 1681708930
transform 1 0 1268 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2104
timestamp 1681708930
transform 1 0 1316 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2105
timestamp 1681708930
transform 1 0 1324 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1893
timestamp 1681708930
transform 1 0 1380 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1920
timestamp 1681708930
transform 1 0 1372 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_2037
timestamp 1681708930
transform 1 0 1372 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2038
timestamp 1681708930
transform 1 0 1380 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_1973
timestamp 1681708930
transform 1 0 1340 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_2039
timestamp 1681708930
transform 1 0 1404 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_1940
timestamp 1681708930
transform 1 0 1412 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_2106
timestamp 1681708930
transform 1 0 1388 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2107
timestamp 1681708930
transform 1 0 1412 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1974
timestamp 1681708930
transform 1 0 1388 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1975
timestamp 1681708930
transform 1 0 1404 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_2152
timestamp 1681708930
transform 1 0 1412 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_1921
timestamp 1681708930
transform 1 0 1444 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_2040
timestamp 1681708930
transform 1 0 1436 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2108
timestamp 1681708930
transform 1 0 1444 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2005
timestamp 1681708930
transform 1 0 1436 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1894
timestamp 1681708930
transform 1 0 1460 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_2007
timestamp 1681708930
transform 1 0 1460 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2041
timestamp 1681708930
transform 1 0 1460 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2008
timestamp 1681708930
transform 1 0 1468 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_1895
timestamp 1681708930
transform 1 0 1508 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_2042
timestamp 1681708930
transform 1 0 1492 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2043
timestamp 1681708930
transform 1 0 1500 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2109
timestamp 1681708930
transform 1 0 1484 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1976
timestamp 1681708930
transform 1 0 1484 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_2110
timestamp 1681708930
transform 1 0 1508 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2111
timestamp 1681708930
transform 1 0 1516 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2021
timestamp 1681708930
transform 1 0 1516 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1922
timestamp 1681708930
transform 1 0 1532 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_2044
timestamp 1681708930
transform 1 0 1532 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2045
timestamp 1681708930
transform 1 0 1564 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_1923
timestamp 1681708930
transform 1 0 1620 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_2046
timestamp 1681708930
transform 1 0 1588 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_1941
timestamp 1681708930
transform 1 0 1596 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_2047
timestamp 1681708930
transform 1 0 1604 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2048
timestamp 1681708930
transform 1 0 1620 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2112
timestamp 1681708930
transform 1 0 1556 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2113
timestamp 1681708930
transform 1 0 1572 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2114
timestamp 1681708930
transform 1 0 1596 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2115
timestamp 1681708930
transform 1 0 1612 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2116
timestamp 1681708930
transform 1 0 1620 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1977
timestamp 1681708930
transform 1 0 1572 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1978
timestamp 1681708930
transform 1 0 1588 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1979
timestamp 1681708930
transform 1 0 1620 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2006
timestamp 1681708930
transform 1 0 1564 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2028
timestamp 1681708930
transform 1 0 1548 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_2022
timestamp 1681708930
transform 1 0 1604 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2029
timestamp 1681708930
transform 1 0 1612 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_2153
timestamp 1681708930
transform 1 0 1636 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2007
timestamp 1681708930
transform 1 0 1636 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_2049
timestamp 1681708930
transform 1 0 1652 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2050
timestamp 1681708930
transform 1 0 1660 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_1954
timestamp 1681708930
transform 1 0 1660 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1881
timestamp 1681708930
transform 1 0 1724 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1924
timestamp 1681708930
transform 1 0 1756 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1942
timestamp 1681708930
transform 1 0 1676 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_2051
timestamp 1681708930
transform 1 0 1756 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_1943
timestamp 1681708930
transform 1 0 1780 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_2052
timestamp 1681708930
transform 1 0 1796 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2053
timestamp 1681708930
transform 1 0 1804 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2054
timestamp 1681708930
transform 1 0 1820 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2055
timestamp 1681708930
transform 1 0 1828 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2117
timestamp 1681708930
transform 1 0 1668 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2118
timestamp 1681708930
transform 1 0 1676 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2119
timestamp 1681708930
transform 1 0 1732 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2120
timestamp 1681708930
transform 1 0 1772 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2121
timestamp 1681708930
transform 1 0 1780 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1955
timestamp 1681708930
transform 1 0 1788 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1980
timestamp 1681708930
transform 1 0 1668 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1981
timestamp 1681708930
transform 1 0 1732 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1982
timestamp 1681708930
transform 1 0 1772 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1956
timestamp 1681708930
transform 1 0 1804 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_2122
timestamp 1681708930
transform 1 0 1812 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1957
timestamp 1681708930
transform 1 0 1828 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1983
timestamp 1681708930
transform 1 0 1820 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1896
timestamp 1681708930
transform 1 0 1876 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_2056
timestamp 1681708930
transform 1 0 1860 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_1944
timestamp 1681708930
transform 1 0 1868 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1897
timestamp 1681708930
transform 1 0 1916 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1882
timestamp 1681708930
transform 1 0 2124 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1898
timestamp 1681708930
transform 1 0 2020 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1899
timestamp 1681708930
transform 1 0 2044 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1900
timestamp 1681708930
transform 1 0 2076 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1901
timestamp 1681708930
transform 1 0 2116 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1925
timestamp 1681708930
transform 1 0 1932 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1926
timestamp 1681708930
transform 1 0 1956 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_2057
timestamp 1681708930
transform 1 0 1892 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2058
timestamp 1681708930
transform 1 0 1900 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2123
timestamp 1681708930
transform 1 0 1860 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2124
timestamp 1681708930
transform 1 0 1868 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2125
timestamp 1681708930
transform 1 0 1884 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1958
timestamp 1681708930
transform 1 0 1892 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_2126
timestamp 1681708930
transform 1 0 1900 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1959
timestamp 1681708930
transform 1 0 1908 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_2059
timestamp 1681708930
transform 1 0 1932 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_1945
timestamp 1681708930
transform 1 0 1980 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1946
timestamp 1681708930
transform 1 0 2012 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_2060
timestamp 1681708930
transform 1 0 2020 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2127
timestamp 1681708930
transform 1 0 1916 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2128
timestamp 1681708930
transform 1 0 1956 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1984
timestamp 1681708930
transform 1 0 1892 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1960
timestamp 1681708930
transform 1 0 1996 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1927
timestamp 1681708930
transform 1 0 2084 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1928
timestamp 1681708930
transform 1 0 2116 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1902
timestamp 1681708930
transform 1 0 2156 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_2061
timestamp 1681708930
transform 1 0 2116 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2062
timestamp 1681708930
transform 1 0 2132 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2129
timestamp 1681708930
transform 1 0 2012 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2130
timestamp 1681708930
transform 1 0 2028 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2131
timestamp 1681708930
transform 1 0 2036 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2132
timestamp 1681708930
transform 1 0 2068 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1985
timestamp 1681708930
transform 1 0 1916 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1986
timestamp 1681708930
transform 1 0 1956 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1961
timestamp 1681708930
transform 1 0 2116 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1962
timestamp 1681708930
transform 1 0 2132 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_2063
timestamp 1681708930
transform 1 0 2180 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2064
timestamp 1681708930
transform 1 0 2188 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2133
timestamp 1681708930
transform 1 0 2148 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1987
timestamp 1681708930
transform 1 0 2028 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1988
timestamp 1681708930
transform 1 0 2068 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1989
timestamp 1681708930
transform 1 0 2084 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2008
timestamp 1681708930
transform 1 0 2044 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2009
timestamp 1681708930
transform 1 0 2068 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1883
timestamp 1681708930
transform 1 0 2300 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_2065
timestamp 1681708930
transform 1 0 2212 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2066
timestamp 1681708930
transform 1 0 2300 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2134
timestamp 1681708930
transform 1 0 2196 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1963
timestamp 1681708930
transform 1 0 2212 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_2135
timestamp 1681708930
transform 1 0 2236 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2136
timestamp 1681708930
transform 1 0 2292 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2137
timestamp 1681708930
transform 1 0 2300 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1990
timestamp 1681708930
transform 1 0 2196 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1991
timestamp 1681708930
transform 1 0 2236 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2010
timestamp 1681708930
transform 1 0 2180 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1903
timestamp 1681708930
transform 1 0 2388 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1929
timestamp 1681708930
transform 1 0 2380 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_2009
timestamp 1681708930
transform 1 0 2388 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2067
timestamp 1681708930
transform 1 0 2380 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2154
timestamp 1681708930
transform 1 0 2388 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2011
timestamp 1681708930
transform 1 0 2388 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1930
timestamp 1681708930
transform 1 0 2404 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1931
timestamp 1681708930
transform 1 0 2428 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_2010
timestamp 1681708930
transform 1 0 2444 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2068
timestamp 1681708930
transform 1 0 2436 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_1992
timestamp 1681708930
transform 1 0 2412 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_2155
timestamp 1681708930
transform 1 0 2420 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2163
timestamp 1681708930
transform 1 0 2412 0 1 1305
box -2 -2 2 2
use M3_M2  M3_M2_1904
timestamp 1681708930
transform 1 0 2460 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_2011
timestamp 1681708930
transform 1 0 2460 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_1905
timestamp 1681708930
transform 1 0 2516 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1932
timestamp 1681708930
transform 1 0 2500 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_2069
timestamp 1681708930
transform 1 0 2484 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2070
timestamp 1681708930
transform 1 0 2500 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2071
timestamp 1681708930
transform 1 0 2516 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2138
timestamp 1681708930
transform 1 0 2460 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2139
timestamp 1681708930
transform 1 0 2468 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1964
timestamp 1681708930
transform 1 0 2484 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_2140
timestamp 1681708930
transform 1 0 2500 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1993
timestamp 1681708930
transform 1 0 2468 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1994
timestamp 1681708930
transform 1 0 2500 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1947
timestamp 1681708930
transform 1 0 2548 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_2072
timestamp 1681708930
transform 1 0 2556 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2141
timestamp 1681708930
transform 1 0 2524 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2142
timestamp 1681708930
transform 1 0 2540 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2156
timestamp 1681708930
transform 1 0 2516 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2157
timestamp 1681708930
transform 1 0 2524 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2012
timestamp 1681708930
transform 1 0 2460 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2013
timestamp 1681708930
transform 1 0 2484 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2014
timestamp 1681708930
transform 1 0 2524 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2023
timestamp 1681708930
transform 1 0 2516 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1965
timestamp 1681708930
transform 1 0 2548 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2015
timestamp 1681708930
transform 1 0 2556 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1906
timestamp 1681708930
transform 1 0 2596 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_2073
timestamp 1681708930
transform 1 0 2572 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2074
timestamp 1681708930
transform 1 0 2628 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_1966
timestamp 1681708930
transform 1 0 2572 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_2143
timestamp 1681708930
transform 1 0 2580 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_1967
timestamp 1681708930
transform 1 0 2596 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_2158
timestamp 1681708930
transform 1 0 2572 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_1995
timestamp 1681708930
transform 1 0 2580 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2016
timestamp 1681708930
transform 1 0 2572 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1996
timestamp 1681708930
transform 1 0 2628 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2024
timestamp 1681708930
transform 1 0 2596 0 1 1295
box -3 -3 3 3
use top_mod_new_VIA0  top_mod_new_VIA0_26
timestamp 1681708930
transform 1 0 24 0 1 1270
box -10 -3 10 3
use FILL  FILL_688
timestamp 1681708930
transform 1 0 72 0 -1 1370
box -8 -3 16 105
use FILL  FILL_690
timestamp 1681708930
transform 1 0 80 0 -1 1370
box -8 -3 16 105
use FILL  FILL_692
timestamp 1681708930
transform 1 0 88 0 -1 1370
box -8 -3 16 105
use FILL  FILL_694
timestamp 1681708930
transform 1 0 96 0 -1 1370
box -8 -3 16 105
use FILL  FILL_711
timestamp 1681708930
transform 1 0 104 0 -1 1370
box -8 -3 16 105
use AOI21X1  AOI21X1_30
timestamp 1681708930
transform -1 0 144 0 -1 1370
box -7 -3 39 105
use INVX2  INVX2_123
timestamp 1681708930
transform -1 0 160 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_124
timestamp 1681708930
transform -1 0 176 0 -1 1370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_44
timestamp 1681708930
transform 1 0 176 0 -1 1370
box -8 -3 104 105
use FILL  FILL_712
timestamp 1681708930
transform 1 0 272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_713
timestamp 1681708930
transform 1 0 280 0 -1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_47
timestamp 1681708930
transform 1 0 288 0 -1 1370
box -8 -3 32 105
use NAND3X1  NAND3X1_74
timestamp 1681708930
transform 1 0 312 0 -1 1370
box -8 -3 40 105
use FILL  FILL_714
timestamp 1681708930
transform 1 0 344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_716
timestamp 1681708930
transform 1 0 352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_718
timestamp 1681708930
transform 1 0 360 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_126
timestamp 1681708930
transform 1 0 368 0 -1 1370
box -9 -3 26 105
use FILL  FILL_727
timestamp 1681708930
transform 1 0 384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_728
timestamp 1681708930
transform 1 0 392 0 -1 1370
box -8 -3 16 105
use FILL  FILL_729
timestamp 1681708930
transform 1 0 400 0 -1 1370
box -8 -3 16 105
use XOR2X1  XOR2X1_91
timestamp 1681708930
transform -1 0 464 0 -1 1370
box -8 -3 64 105
use NAND3X1  NAND3X1_76
timestamp 1681708930
transform 1 0 464 0 -1 1370
box -8 -3 40 105
use FILL  FILL_730
timestamp 1681708930
transform 1 0 496 0 -1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_77
timestamp 1681708930
transform -1 0 536 0 -1 1370
box -8 -3 40 105
use FILL  FILL_731
timestamp 1681708930
transform 1 0 536 0 -1 1370
box -8 -3 16 105
use FILL  FILL_732
timestamp 1681708930
transform 1 0 544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_733
timestamp 1681708930
transform 1 0 552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_735
timestamp 1681708930
transform 1 0 560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_737
timestamp 1681708930
transform 1 0 568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_738
timestamp 1681708930
transform 1 0 576 0 -1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_78
timestamp 1681708930
transform -1 0 616 0 -1 1370
box -8 -3 40 105
use FILL  FILL_739
timestamp 1681708930
transform 1 0 616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_740
timestamp 1681708930
transform 1 0 624 0 -1 1370
box -8 -3 16 105
use FILL  FILL_742
timestamp 1681708930
transform 1 0 632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_744
timestamp 1681708930
transform 1 0 640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_745
timestamp 1681708930
transform 1 0 648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_746
timestamp 1681708930
transform 1 0 656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_747
timestamp 1681708930
transform 1 0 664 0 -1 1370
box -8 -3 16 105
use FILL  FILL_748
timestamp 1681708930
transform 1 0 672 0 -1 1370
box -8 -3 16 105
use FILL  FILL_749
timestamp 1681708930
transform 1 0 680 0 -1 1370
box -8 -3 16 105
use FILL  FILL_750
timestamp 1681708930
transform 1 0 688 0 -1 1370
box -8 -3 16 105
use FILL  FILL_751
timestamp 1681708930
transform 1 0 696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_752
timestamp 1681708930
transform 1 0 704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_753
timestamp 1681708930
transform 1 0 712 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_2030
timestamp 1681708930
transform 1 0 732 0 1 1275
box -3 -3 3 3
use FILL  FILL_754
timestamp 1681708930
transform 1 0 720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_755
timestamp 1681708930
transform 1 0 728 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_36
timestamp 1681708930
transform 1 0 736 0 -1 1370
box -8 -3 46 105
use FILL  FILL_805
timestamp 1681708930
transform 1 0 776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_806
timestamp 1681708930
transform 1 0 784 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_46
timestamp 1681708930
transform -1 0 888 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_47
timestamp 1681708930
transform 1 0 888 0 -1 1370
box -8 -3 104 105
use FILL  FILL_807
timestamp 1681708930
transform 1 0 984 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_133
timestamp 1681708930
transform 1 0 992 0 -1 1370
box -9 -3 26 105
use FILL  FILL_808
timestamp 1681708930
transform 1 0 1008 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_37
timestamp 1681708930
transform 1 0 1016 0 -1 1370
box -8 -3 46 105
use M3_M2  M3_M2_2031
timestamp 1681708930
transform 1 0 1068 0 1 1275
box -3 -3 3 3
use FILL  FILL_809
timestamp 1681708930
transform 1 0 1056 0 -1 1370
box -8 -3 16 105
use FILL  FILL_810
timestamp 1681708930
transform 1 0 1064 0 -1 1370
box -8 -3 16 105
use FILL  FILL_811
timestamp 1681708930
transform 1 0 1072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_812
timestamp 1681708930
transform 1 0 1080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_813
timestamp 1681708930
transform 1 0 1088 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_38
timestamp 1681708930
transform 1 0 1096 0 -1 1370
box -8 -3 46 105
use M3_M2  M3_M2_2032
timestamp 1681708930
transform 1 0 1148 0 1 1275
box -3 -3 3 3
use FILL  FILL_814
timestamp 1681708930
transform 1 0 1136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_815
timestamp 1681708930
transform 1 0 1144 0 -1 1370
box -8 -3 16 105
use FILL  FILL_816
timestamp 1681708930
transform 1 0 1152 0 -1 1370
box -8 -3 16 105
use FILL  FILL_817
timestamp 1681708930
transform 1 0 1160 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_39
timestamp 1681708930
transform 1 0 1168 0 -1 1370
box -8 -3 46 105
use FILL  FILL_818
timestamp 1681708930
transform 1 0 1208 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_2033
timestamp 1681708930
transform 1 0 1228 0 1 1275
box -3 -3 3 3
use FILL  FILL_819
timestamp 1681708930
transform 1 0 1216 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_48
timestamp 1681708930
transform 1 0 1224 0 -1 1370
box -8 -3 104 105
use XOR2X1  XOR2X1_97
timestamp 1681708930
transform -1 0 1376 0 -1 1370
box -8 -3 64 105
use OAI21X1  OAI21X1_56
timestamp 1681708930
transform 1 0 1376 0 -1 1370
box -8 -3 34 105
use NAND2X1  NAND2X1_50
timestamp 1681708930
transform -1 0 1432 0 -1 1370
box -8 -3 32 105
use FILL  FILL_820
timestamp 1681708930
transform 1 0 1432 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_134
timestamp 1681708930
transform 1 0 1440 0 -1 1370
box -9 -3 26 105
use FILL  FILL_821
timestamp 1681708930
transform 1 0 1456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_822
timestamp 1681708930
transform 1 0 1464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_823
timestamp 1681708930
transform 1 0 1472 0 -1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_49
timestamp 1681708930
transform 1 0 1480 0 -1 1370
box -8 -3 32 105
use INVX2  INVX2_135
timestamp 1681708930
transform -1 0 1520 0 -1 1370
box -9 -3 26 105
use FILL  FILL_824
timestamp 1681708930
transform 1 0 1520 0 -1 1370
box -8 -3 16 105
use FILL  FILL_825
timestamp 1681708930
transform 1 0 1528 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_40
timestamp 1681708930
transform 1 0 1536 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_41
timestamp 1681708930
transform -1 0 1616 0 -1 1370
box -8 -3 46 105
use NAND2X1  NAND2X1_51
timestamp 1681708930
transform 1 0 1616 0 -1 1370
box -8 -3 32 105
use INVX2  INVX2_136
timestamp 1681708930
transform -1 0 1656 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_137
timestamp 1681708930
transform 1 0 1656 0 -1 1370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_49
timestamp 1681708930
transform -1 0 1768 0 -1 1370
box -8 -3 104 105
use INVX2  INVX2_138
timestamp 1681708930
transform -1 0 1784 0 -1 1370
box -9 -3 26 105
use FILL  FILL_826
timestamp 1681708930
transform 1 0 1784 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_42
timestamp 1681708930
transform -1 0 1832 0 -1 1370
box -8 -3 46 105
use FILL  FILL_827
timestamp 1681708930
transform 1 0 1832 0 -1 1370
box -8 -3 16 105
use FILL  FILL_829
timestamp 1681708930
transform 1 0 1840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_831
timestamp 1681708930
transform 1 0 1848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_868
timestamp 1681708930
transform 1 0 1856 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_2034
timestamp 1681708930
transform 1 0 1908 0 1 1275
box -3 -3 3 3
use AOI22X1  AOI22X1_45
timestamp 1681708930
transform -1 0 1904 0 -1 1370
box -8 -3 46 105
use INVX2  INVX2_143
timestamp 1681708930
transform 1 0 1904 0 -1 1370
box -9 -3 26 105
use M3_M2  M3_M2_2035
timestamp 1681708930
transform 1 0 2020 0 1 1275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_51
timestamp 1681708930
transform 1 0 1920 0 -1 1370
box -8 -3 104 105
use INVX2  INVX2_144
timestamp 1681708930
transform 1 0 2016 0 -1 1370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_52
timestamp 1681708930
transform -1 0 2128 0 -1 1370
box -8 -3 104 105
use M3_M2  M3_M2_2036
timestamp 1681708930
transform 1 0 2148 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2037
timestamp 1681708930
transform 1 0 2180 0 1 1275
box -3 -3 3 3
use XNOR2X1  XNOR2X1_33
timestamp 1681708930
transform -1 0 2184 0 -1 1370
box -8 -3 64 105
use INVX2  INVX2_145
timestamp 1681708930
transform 1 0 2184 0 -1 1370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_53
timestamp 1681708930
transform 1 0 2200 0 -1 1370
box -8 -3 104 105
use XNOR2X1  XNOR2X1_34
timestamp 1681708930
transform -1 0 2352 0 -1 1370
box -8 -3 64 105
use OR2X1  OR2X1_12
timestamp 1681708930
transform -1 0 2384 0 -1 1370
box -8 -3 40 105
use FILL  FILL_869
timestamp 1681708930
transform 1 0 2384 0 -1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_82
timestamp 1681708930
transform -1 0 2424 0 -1 1370
box -8 -3 40 105
use INVX2  INVX2_146
timestamp 1681708930
transform -1 0 2440 0 -1 1370
box -9 -3 26 105
use NOR2X1  NOR2X1_50
timestamp 1681708930
transform 1 0 2440 0 -1 1370
box -8 -3 32 105
use AOI21X1  AOI21X1_33
timestamp 1681708930
transform -1 0 2496 0 -1 1370
box -7 -3 39 105
use NAND2X1  NAND2X1_53
timestamp 1681708930
transform 1 0 2496 0 -1 1370
box -8 -3 32 105
use OAI21X1  OAI21X1_58
timestamp 1681708930
transform -1 0 2552 0 -1 1370
box -8 -3 34 105
use NAND2X1  NAND2X1_54
timestamp 1681708930
transform 1 0 2552 0 -1 1370
box -8 -3 32 105
use XNOR2X1  XNOR2X1_35
timestamp 1681708930
transform -1 0 2632 0 -1 1370
box -8 -3 64 105
use FILL  FILL_870
timestamp 1681708930
transform 1 0 2632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_872
timestamp 1681708930
transform 1 0 2640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_874
timestamp 1681708930
transform 1 0 2648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_876
timestamp 1681708930
transform 1 0 2656 0 -1 1370
box -8 -3 16 105
use top_mod_new_VIA0  top_mod_new_VIA0_27
timestamp 1681708930
transform 1 0 2712 0 1 1270
box -10 -3 10 3
use M2_M1  M2_M1_2164
timestamp 1681708930
transform 1 0 132 0 1 1235
box -2 -2 2 2
use M3_M2  M3_M2_2094
timestamp 1681708930
transform 1 0 116 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2180
timestamp 1681708930
transform 1 0 116 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2249
timestamp 1681708930
transform 1 0 108 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2072
timestamp 1681708930
transform 1 0 172 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2073
timestamp 1681708930
transform 1 0 188 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_2168
timestamp 1681708930
transform 1 0 140 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_2095
timestamp 1681708930
transform 1 0 148 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2169
timestamp 1681708930
transform 1 0 156 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_2096
timestamp 1681708930
transform 1 0 164 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2181
timestamp 1681708930
transform 1 0 140 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2155
timestamp 1681708930
transform 1 0 132 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2129
timestamp 1681708930
transform 1 0 156 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_2182
timestamp 1681708930
transform 1 0 164 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2250
timestamp 1681708930
transform 1 0 164 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2156
timestamp 1681708930
transform 1 0 164 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_2170
timestamp 1681708930
transform 1 0 188 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_2130
timestamp 1681708930
transform 1 0 188 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_2183
timestamp 1681708930
transform 1 0 228 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2184
timestamp 1681708930
transform 1 0 284 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2185
timestamp 1681708930
transform 1 0 300 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2251
timestamp 1681708930
transform 1 0 188 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2252
timestamp 1681708930
transform 1 0 204 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2253
timestamp 1681708930
transform 1 0 292 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2157
timestamp 1681708930
transform 1 0 188 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2158
timestamp 1681708930
transform 1 0 204 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2159
timestamp 1681708930
transform 1 0 268 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_2171
timestamp 1681708930
transform 1 0 332 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2186
timestamp 1681708930
transform 1 0 324 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2187
timestamp 1681708930
transform 1 0 332 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2160
timestamp 1681708930
transform 1 0 324 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2182
timestamp 1681708930
transform 1 0 324 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_2254
timestamp 1681708930
transform 1 0 348 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2161
timestamp 1681708930
transform 1 0 348 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_2255
timestamp 1681708930
transform 1 0 372 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2162
timestamp 1681708930
transform 1 0 364 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2183
timestamp 1681708930
transform 1 0 356 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_2188
timestamp 1681708930
transform 1 0 412 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2256
timestamp 1681708930
transform 1 0 420 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2074
timestamp 1681708930
transform 1 0 436 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2075
timestamp 1681708930
transform 1 0 452 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2076
timestamp 1681708930
transform 1 0 468 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_2172
timestamp 1681708930
transform 1 0 436 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2173
timestamp 1681708930
transform 1 0 468 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2189
timestamp 1681708930
transform 1 0 436 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2190
timestamp 1681708930
transform 1 0 452 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2257
timestamp 1681708930
transform 1 0 444 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2163
timestamp 1681708930
transform 1 0 436 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_2258
timestamp 1681708930
transform 1 0 468 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2259
timestamp 1681708930
transform 1 0 476 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2164
timestamp 1681708930
transform 1 0 476 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2184
timestamp 1681708930
transform 1 0 452 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2038
timestamp 1681708930
transform 1 0 492 0 1 1265
box -3 -3 3 3
use M2_M1  M2_M1_2260
timestamp 1681708930
transform 1 0 492 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2097
timestamp 1681708930
transform 1 0 516 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2077
timestamp 1681708930
transform 1 0 540 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2078
timestamp 1681708930
transform 1 0 572 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2098
timestamp 1681708930
transform 1 0 556 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2191
timestamp 1681708930
transform 1 0 516 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2192
timestamp 1681708930
transform 1 0 524 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2193
timestamp 1681708930
transform 1 0 540 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2194
timestamp 1681708930
transform 1 0 556 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2185
timestamp 1681708930
transform 1 0 508 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2131
timestamp 1681708930
transform 1 0 564 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_2195
timestamp 1681708930
transform 1 0 580 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2196
timestamp 1681708930
transform 1 0 604 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2261
timestamp 1681708930
transform 1 0 564 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2262
timestamp 1681708930
transform 1 0 572 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2141
timestamp 1681708930
transform 1 0 580 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_2263
timestamp 1681708930
transform 1 0 588 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2264
timestamp 1681708930
transform 1 0 596 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2142
timestamp 1681708930
transform 1 0 604 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2079
timestamp 1681708930
transform 1 0 652 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_2174
timestamp 1681708930
transform 1 0 652 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2197
timestamp 1681708930
transform 1 0 644 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2198
timestamp 1681708930
transform 1 0 652 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2265
timestamp 1681708930
transform 1 0 620 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2165
timestamp 1681708930
transform 1 0 564 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2143
timestamp 1681708930
transform 1 0 628 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_2266
timestamp 1681708930
transform 1 0 636 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2166
timestamp 1681708930
transform 1 0 620 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_2267
timestamp 1681708930
transform 1 0 660 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2311
timestamp 1681708930
transform 1 0 628 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_2186
timestamp 1681708930
transform 1 0 620 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2167
timestamp 1681708930
transform 1 0 644 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2039
timestamp 1681708930
transform 1 0 732 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2132
timestamp 1681708930
transform 1 0 724 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2040
timestamp 1681708930
transform 1 0 804 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2047
timestamp 1681708930
transform 1 0 772 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2048
timestamp 1681708930
transform 1 0 788 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2049
timestamp 1681708930
transform 1 0 836 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2061
timestamp 1681708930
transform 1 0 804 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2062
timestamp 1681708930
transform 1 0 844 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2080
timestamp 1681708930
transform 1 0 844 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2099
timestamp 1681708930
transform 1 0 756 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2100
timestamp 1681708930
transform 1 0 796 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2199
timestamp 1681708930
transform 1 0 740 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2200
timestamp 1681708930
transform 1 0 756 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2201
timestamp 1681708930
transform 1 0 764 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2202
timestamp 1681708930
transform 1 0 796 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2268
timestamp 1681708930
transform 1 0 708 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2269
timestamp 1681708930
transform 1 0 724 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2168
timestamp 1681708930
transform 1 0 708 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_2312
timestamp 1681708930
transform 1 0 716 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_2187
timestamp 1681708930
transform 1 0 708 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2144
timestamp 1681708930
transform 1 0 740 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_2270
timestamp 1681708930
transform 1 0 748 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2145
timestamp 1681708930
transform 1 0 804 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2063
timestamp 1681708930
transform 1 0 876 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2050
timestamp 1681708930
transform 1 0 948 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2081
timestamp 1681708930
transform 1 0 876 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2082
timestamp 1681708930
transform 1 0 916 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2101
timestamp 1681708930
transform 1 0 884 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2102
timestamp 1681708930
transform 1 0 908 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2103
timestamp 1681708930
transform 1 0 940 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2203
timestamp 1681708930
transform 1 0 884 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2204
timestamp 1681708930
transform 1 0 916 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2205
timestamp 1681708930
transform 1 0 940 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2271
timestamp 1681708930
transform 1 0 844 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2272
timestamp 1681708930
transform 1 0 860 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2169
timestamp 1681708930
transform 1 0 820 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2188
timestamp 1681708930
transform 1 0 740 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2189
timestamp 1681708930
transform 1 0 764 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2190
timestamp 1681708930
transform 1 0 852 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2191
timestamp 1681708930
transform 1 0 884 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2133
timestamp 1681708930
transform 1 0 948 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2041
timestamp 1681708930
transform 1 0 1020 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2051
timestamp 1681708930
transform 1 0 980 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2052
timestamp 1681708930
transform 1 0 1028 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2053
timestamp 1681708930
transform 1 0 1052 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2064
timestamp 1681708930
transform 1 0 980 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2054
timestamp 1681708930
transform 1 0 1092 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2083
timestamp 1681708930
transform 1 0 1092 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2104
timestamp 1681708930
transform 1 0 1084 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2206
timestamp 1681708930
transform 1 0 964 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2207
timestamp 1681708930
transform 1 0 1004 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2208
timestamp 1681708930
transform 1 0 1060 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2134
timestamp 1681708930
transform 1 0 1068 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2042
timestamp 1681708930
transform 1 0 1164 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2043
timestamp 1681708930
transform 1 0 1188 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2044
timestamp 1681708930
transform 1 0 1236 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2055
timestamp 1681708930
transform 1 0 1188 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2065
timestamp 1681708930
transform 1 0 1148 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2105
timestamp 1681708930
transform 1 0 1132 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2106
timestamp 1681708930
transform 1 0 1172 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2056
timestamp 1681708930
transform 1 0 1316 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2066
timestamp 1681708930
transform 1 0 1244 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2067
timestamp 1681708930
transform 1 0 1260 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2084
timestamp 1681708930
transform 1 0 1292 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2085
timestamp 1681708930
transform 1 0 1348 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2107
timestamp 1681708930
transform 1 0 1244 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2108
timestamp 1681708930
transform 1 0 1284 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2109
timestamp 1681708930
transform 1 0 1332 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2209
timestamp 1681708930
transform 1 0 1092 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2210
timestamp 1681708930
transform 1 0 1100 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2211
timestamp 1681708930
transform 1 0 1124 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2212
timestamp 1681708930
transform 1 0 1132 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2213
timestamp 1681708930
transform 1 0 1172 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2214
timestamp 1681708930
transform 1 0 1228 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2215
timestamp 1681708930
transform 1 0 1236 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2216
timestamp 1681708930
transform 1 0 1244 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2217
timestamp 1681708930
transform 1 0 1284 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2218
timestamp 1681708930
transform 1 0 1340 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2219
timestamp 1681708930
transform 1 0 1348 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2146
timestamp 1681708930
transform 1 0 964 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_2273
timestamp 1681708930
transform 1 0 980 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2147
timestamp 1681708930
transform 1 0 1012 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_2274
timestamp 1681708930
transform 1 0 1068 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2170
timestamp 1681708930
transform 1 0 1012 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_2275
timestamp 1681708930
transform 1 0 1116 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2148
timestamp 1681708930
transform 1 0 1124 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2192
timestamp 1681708930
transform 1 0 1068 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2193
timestamp 1681708930
transform 1 0 1092 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2194
timestamp 1681708930
transform 1 0 1108 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_2276
timestamp 1681708930
transform 1 0 1148 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2171
timestamp 1681708930
transform 1 0 1220 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_2277
timestamp 1681708930
transform 1 0 1260 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2278
timestamp 1681708930
transform 1 0 1348 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2172
timestamp 1681708930
transform 1 0 1348 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2086
timestamp 1681708930
transform 1 0 1428 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2110
timestamp 1681708930
transform 1 0 1428 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2220
timestamp 1681708930
transform 1 0 1428 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2221
timestamp 1681708930
transform 1 0 1436 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2279
timestamp 1681708930
transform 1 0 1396 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2280
timestamp 1681708930
transform 1 0 1404 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2195
timestamp 1681708930
transform 1 0 1380 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_2165
timestamp 1681708930
transform 1 0 1460 0 1 1235
box -2 -2 2 2
use M3_M2  M3_M2_2111
timestamp 1681708930
transform 1 0 1460 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2087
timestamp 1681708930
transform 1 0 1484 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_2175
timestamp 1681708930
transform 1 0 1468 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2248
timestamp 1681708930
transform 1 0 1460 0 1 1214
box -2 -2 2 2
use M2_M1  M2_M1_2281
timestamp 1681708930
transform 1 0 1460 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2176
timestamp 1681708930
transform 1 0 1500 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2313
timestamp 1681708930
transform 1 0 1532 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2282
timestamp 1681708930
transform 1 0 1548 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2112
timestamp 1681708930
transform 1 0 1564 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2314
timestamp 1681708930
transform 1 0 1564 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2283
timestamp 1681708930
transform 1 0 1620 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2057
timestamp 1681708930
transform 1 0 1740 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2113
timestamp 1681708930
transform 1 0 1692 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2114
timestamp 1681708930
transform 1 0 1732 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2222
timestamp 1681708930
transform 1 0 1636 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2223
timestamp 1681708930
transform 1 0 1692 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2224
timestamp 1681708930
transform 1 0 1732 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2149
timestamp 1681708930
transform 1 0 1636 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_2284
timestamp 1681708930
transform 1 0 1716 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2315
timestamp 1681708930
transform 1 0 1628 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2225
timestamp 1681708930
transform 1 0 1748 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2150
timestamp 1681708930
transform 1 0 1748 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2196
timestamp 1681708930
transform 1 0 1740 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2045
timestamp 1681708930
transform 1 0 1796 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2046
timestamp 1681708930
transform 1 0 1820 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2088
timestamp 1681708930
transform 1 0 1780 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2089
timestamp 1681708930
transform 1 0 1804 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2115
timestamp 1681708930
transform 1 0 1812 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2116
timestamp 1681708930
transform 1 0 1836 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2117
timestamp 1681708930
transform 1 0 1860 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2226
timestamp 1681708930
transform 1 0 1788 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2227
timestamp 1681708930
transform 1 0 1812 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2228
timestamp 1681708930
transform 1 0 1836 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2229
timestamp 1681708930
transform 1 0 1860 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2285
timestamp 1681708930
transform 1 0 1772 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2286
timestamp 1681708930
transform 1 0 1780 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2287
timestamp 1681708930
transform 1 0 1796 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2288
timestamp 1681708930
transform 1 0 1812 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2197
timestamp 1681708930
transform 1 0 1812 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_2230
timestamp 1681708930
transform 1 0 1876 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2118
timestamp 1681708930
transform 1 0 1932 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2090
timestamp 1681708930
transform 1 0 1988 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_2231
timestamp 1681708930
transform 1 0 1900 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2232
timestamp 1681708930
transform 1 0 1932 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2289
timestamp 1681708930
transform 1 0 1884 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2173
timestamp 1681708930
transform 1 0 1884 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2198
timestamp 1681708930
transform 1 0 1876 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2135
timestamp 1681708930
transform 1 0 1940 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2136
timestamp 1681708930
transform 1 0 1964 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_2290
timestamp 1681708930
transform 1 0 1932 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2291
timestamp 1681708930
transform 1 0 1940 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2174
timestamp 1681708930
transform 1 0 1932 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2199
timestamp 1681708930
transform 1 0 1900 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2200
timestamp 1681708930
transform 1 0 1964 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_2233
timestamp 1681708930
transform 1 0 1996 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2201
timestamp 1681708930
transform 1 0 1996 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_2234
timestamp 1681708930
transform 1 0 2028 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2235
timestamp 1681708930
transform 1 0 2044 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2292
timestamp 1681708930
transform 1 0 2012 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2293
timestamp 1681708930
transform 1 0 2020 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2151
timestamp 1681708930
transform 1 0 2028 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2202
timestamp 1681708930
transform 1 0 2020 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2137
timestamp 1681708930
transform 1 0 2060 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_2294
timestamp 1681708930
transform 1 0 2060 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2203
timestamp 1681708930
transform 1 0 2052 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2091
timestamp 1681708930
transform 1 0 2076 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2119
timestamp 1681708930
transform 1 0 2092 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2236
timestamp 1681708930
transform 1 0 2092 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2120
timestamp 1681708930
transform 1 0 2124 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2068
timestamp 1681708930
transform 1 0 2140 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2121
timestamp 1681708930
transform 1 0 2156 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2237
timestamp 1681708930
transform 1 0 2140 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2138
timestamp 1681708930
transform 1 0 2148 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_2238
timestamp 1681708930
transform 1 0 2156 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2295
timestamp 1681708930
transform 1 0 2140 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2296
timestamp 1681708930
transform 1 0 2148 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2152
timestamp 1681708930
transform 1 0 2156 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_2297
timestamp 1681708930
transform 1 0 2164 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2204
timestamp 1681708930
transform 1 0 2140 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2122
timestamp 1681708930
transform 1 0 2188 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2239
timestamp 1681708930
transform 1 0 2236 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2139
timestamp 1681708930
transform 1 0 2276 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2069
timestamp 1681708930
transform 1 0 2292 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_2240
timestamp 1681708930
transform 1 0 2284 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2298
timestamp 1681708930
transform 1 0 2276 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2299
timestamp 1681708930
transform 1 0 2332 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2300
timestamp 1681708930
transform 1 0 2340 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2205
timestamp 1681708930
transform 1 0 2332 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2123
timestamp 1681708930
transform 1 0 2356 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2241
timestamp 1681708930
transform 1 0 2348 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2140
timestamp 1681708930
transform 1 0 2364 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_2301
timestamp 1681708930
transform 1 0 2356 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2175
timestamp 1681708930
transform 1 0 2348 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2070
timestamp 1681708930
transform 1 0 2396 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2071
timestamp 1681708930
transform 1 0 2412 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2092
timestamp 1681708930
transform 1 0 2396 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2124
timestamp 1681708930
transform 1 0 2388 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2177
timestamp 1681708930
transform 1 0 2396 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2302
timestamp 1681708930
transform 1 0 2380 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2058
timestamp 1681708930
transform 1 0 2436 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2059
timestamp 1681708930
transform 1 0 2452 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2125
timestamp 1681708930
transform 1 0 2428 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2242
timestamp 1681708930
transform 1 0 2428 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2093
timestamp 1681708930
transform 1 0 2444 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2126
timestamp 1681708930
transform 1 0 2452 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2243
timestamp 1681708930
transform 1 0 2452 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2244
timestamp 1681708930
transform 1 0 2476 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2303
timestamp 1681708930
transform 1 0 2428 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2304
timestamp 1681708930
transform 1 0 2436 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2305
timestamp 1681708930
transform 1 0 2444 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2306
timestamp 1681708930
transform 1 0 2468 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2176
timestamp 1681708930
transform 1 0 2436 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2153
timestamp 1681708930
transform 1 0 2476 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_2307
timestamp 1681708930
transform 1 0 2484 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2177
timestamp 1681708930
transform 1 0 2484 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2127
timestamp 1681708930
transform 1 0 2500 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2154
timestamp 1681708930
transform 1 0 2500 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2060
timestamp 1681708930
transform 1 0 2540 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_2166
timestamp 1681708930
transform 1 0 2532 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_2167
timestamp 1681708930
transform 1 0 2548 0 1 1235
box -2 -2 2 2
use M3_M2  M3_M2_2128
timestamp 1681708930
transform 1 0 2524 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_2178
timestamp 1681708930
transform 1 0 2532 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2179
timestamp 1681708930
transform 1 0 2556 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2245
timestamp 1681708930
transform 1 0 2540 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2308
timestamp 1681708930
transform 1 0 2516 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2309
timestamp 1681708930
transform 1 0 2524 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2316
timestamp 1681708930
transform 1 0 2500 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_2178
timestamp 1681708930
transform 1 0 2508 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2179
timestamp 1681708930
transform 1 0 2524 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2180
timestamp 1681708930
transform 1 0 2548 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_2246
timestamp 1681708930
transform 1 0 2564 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2181
timestamp 1681708930
transform 1 0 2564 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_2310
timestamp 1681708930
transform 1 0 2596 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2317
timestamp 1681708930
transform 1 0 2580 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2247
timestamp 1681708930
transform 1 0 2620 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2318
timestamp 1681708930
transform 1 0 2652 0 1 1195
box -2 -2 2 2
use top_mod_new_VIA0  top_mod_new_VIA0_28
timestamp 1681708930
transform 1 0 48 0 1 1170
box -10 -3 10 3
use FILL  FILL_877
timestamp 1681708930
transform 1 0 72 0 1 1170
box -8 -3 16 105
use FILL  FILL_878
timestamp 1681708930
transform 1 0 80 0 1 1170
box -8 -3 16 105
use FILL  FILL_879
timestamp 1681708930
transform 1 0 88 0 1 1170
box -8 -3 16 105
use FILL  FILL_880
timestamp 1681708930
transform 1 0 96 0 1 1170
box -8 -3 16 105
use FILL  FILL_881
timestamp 1681708930
transform 1 0 104 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_147
timestamp 1681708930
transform 1 0 112 0 1 1170
box -9 -3 26 105
use NAND3X1  NAND3X1_83
timestamp 1681708930
transform 1 0 128 0 1 1170
box -8 -3 40 105
use OAI21X1  OAI21X1_59
timestamp 1681708930
transform 1 0 160 0 1 1170
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_54
timestamp 1681708930
transform 1 0 192 0 1 1170
box -8 -3 104 105
use AND2X2  AND2X2_2
timestamp 1681708930
transform 1 0 288 0 1 1170
box -8 -3 40 105
use FILL  FILL_882
timestamp 1681708930
transform 1 0 320 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_2206
timestamp 1681708930
transform 1 0 356 0 1 1175
box -3 -3 3 3
use NAND2X1  NAND2X1_55
timestamp 1681708930
transform -1 0 352 0 1 1170
box -8 -3 32 105
use FILL  FILL_883
timestamp 1681708930
transform 1 0 352 0 1 1170
box -8 -3 16 105
use OR2X1  OR2X1_13
timestamp 1681708930
transform 1 0 360 0 1 1170
box -8 -3 40 105
use FILL  FILL_884
timestamp 1681708930
transform 1 0 392 0 1 1170
box -8 -3 16 105
use FILL  FILL_885
timestamp 1681708930
transform 1 0 400 0 1 1170
box -8 -3 16 105
use FILL  FILL_886
timestamp 1681708930
transform 1 0 408 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_2207
timestamp 1681708930
transform 1 0 428 0 1 1175
box -3 -3 3 3
use NAND2X1  NAND2X1_56
timestamp 1681708930
transform 1 0 416 0 1 1170
box -8 -3 32 105
use OAI21X1  OAI21X1_60
timestamp 1681708930
transform 1 0 440 0 1 1170
box -8 -3 34 105
use INVX2  INVX2_148
timestamp 1681708930
transform 1 0 472 0 1 1170
box -9 -3 26 105
use FILL  FILL_887
timestamp 1681708930
transform 1 0 488 0 1 1170
box -8 -3 16 105
use FILL  FILL_888
timestamp 1681708930
transform 1 0 496 0 1 1170
box -8 -3 16 105
use FILL  FILL_889
timestamp 1681708930
transform 1 0 504 0 1 1170
box -8 -3 16 105
use FILL  FILL_890
timestamp 1681708930
transform 1 0 512 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_2208
timestamp 1681708930
transform 1 0 532 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2209
timestamp 1681708930
transform 1 0 556 0 1 1175
box -3 -3 3 3
use AOI22X1  AOI22X1_46
timestamp 1681708930
transform 1 0 520 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_47
timestamp 1681708930
transform -1 0 600 0 1 1170
box -8 -3 46 105
use OR2X1  OR2X1_14
timestamp 1681708930
transform -1 0 632 0 1 1170
box -8 -3 40 105
use NAND2X1  NAND2X1_57
timestamp 1681708930
transform 1 0 632 0 1 1170
box -8 -3 32 105
use M3_M2  M3_M2_2210
timestamp 1681708930
transform 1 0 684 0 1 1175
box -3 -3 3 3
use XOR2X1  XOR2X1_101
timestamp 1681708930
transform -1 0 712 0 1 1170
box -8 -3 64 105
use OR2X1  OR2X1_15
timestamp 1681708930
transform 1 0 712 0 1 1170
box -8 -3 40 105
use INVX2  INVX2_149
timestamp 1681708930
transform 1 0 744 0 1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_55
timestamp 1681708930
transform -1 0 856 0 1 1170
box -8 -3 104 105
use M3_M2  M3_M2_2211
timestamp 1681708930
transform 1 0 908 0 1 1175
box -3 -3 3 3
use XOR2X1  XOR2X1_102
timestamp 1681708930
transform -1 0 912 0 1 1170
box -8 -3 64 105
use M3_M2  M3_M2_2212
timestamp 1681708930
transform 1 0 956 0 1 1175
box -3 -3 3 3
use XOR2X1  XOR2X1_103
timestamp 1681708930
transform 1 0 912 0 1 1170
box -8 -3 64 105
use M3_M2  M3_M2_2213
timestamp 1681708930
transform 1 0 1020 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2214
timestamp 1681708930
transform 1 0 1068 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_56
timestamp 1681708930
transform 1 0 968 0 1 1170
box -8 -3 104 105
use XOR2X1  XOR2X1_104
timestamp 1681708930
transform 1 0 1064 0 1 1170
box -8 -3 64 105
use INVX2  INVX2_150
timestamp 1681708930
transform 1 0 1120 0 1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_57
timestamp 1681708930
transform 1 0 1136 0 1 1170
box -8 -3 104 105
use INVX2  INVX2_151
timestamp 1681708930
transform 1 0 1232 0 1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_58
timestamp 1681708930
transform 1 0 1248 0 1 1170
box -8 -3 104 105
use XOR2X1  XOR2X1_105
timestamp 1681708930
transform -1 0 1400 0 1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_106
timestamp 1681708930
transform 1 0 1400 0 1 1170
box -8 -3 64 105
use FILL  FILL_891
timestamp 1681708930
transform 1 0 1456 0 1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_85
timestamp 1681708930
transform 1 0 1464 0 1 1170
box -8 -3 40 105
use FILL  FILL_944
timestamp 1681708930
transform 1 0 1496 0 1 1170
box -8 -3 16 105
use FILL  FILL_945
timestamp 1681708930
transform 1 0 1504 0 1 1170
box -8 -3 16 105
use FILL  FILL_948
timestamp 1681708930
transform 1 0 1512 0 1 1170
box -8 -3 16 105
use FILL  FILL_950
timestamp 1681708930
transform 1 0 1520 0 1 1170
box -8 -3 16 105
use FILL  FILL_951
timestamp 1681708930
transform 1 0 1528 0 1 1170
box -8 -3 16 105
use FILL  FILL_952
timestamp 1681708930
transform 1 0 1536 0 1 1170
box -8 -3 16 105
use FILL  FILL_953
timestamp 1681708930
transform 1 0 1544 0 1 1170
box -8 -3 16 105
use FILL  FILL_954
timestamp 1681708930
transform 1 0 1552 0 1 1170
box -8 -3 16 105
use FILL  FILL_955
timestamp 1681708930
transform 1 0 1560 0 1 1170
box -8 -3 16 105
use FILL  FILL_956
timestamp 1681708930
transform 1 0 1568 0 1 1170
box -8 -3 16 105
use FILL  FILL_957
timestamp 1681708930
transform 1 0 1576 0 1 1170
box -8 -3 16 105
use FILL  FILL_958
timestamp 1681708930
transform 1 0 1584 0 1 1170
box -8 -3 16 105
use OR2X1  OR2X1_16
timestamp 1681708930
transform -1 0 1624 0 1 1170
box -8 -3 40 105
use FILL  FILL_959
timestamp 1681708930
transform 1 0 1624 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_62
timestamp 1681708930
transform -1 0 1728 0 1 1170
box -8 -3 104 105
use INVX2  INVX2_158
timestamp 1681708930
transform -1 0 1744 0 1 1170
box -9 -3 26 105
use FILL  FILL_960
timestamp 1681708930
transform 1 0 1744 0 1 1170
box -8 -3 16 105
use FILL  FILL_961
timestamp 1681708930
transform 1 0 1752 0 1 1170
box -8 -3 16 105
use FILL  FILL_962
timestamp 1681708930
transform 1 0 1760 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_49
timestamp 1681708930
transform -1 0 1808 0 1 1170
box -8 -3 46 105
use XOR2X1  XOR2X1_112
timestamp 1681708930
transform 1 0 1808 0 1 1170
box -8 -3 64 105
use FILL  FILL_963
timestamp 1681708930
transform 1 0 1864 0 1 1170
box -8 -3 16 105
use FILL  FILL_964
timestamp 1681708930
transform 1 0 1872 0 1 1170
box -8 -3 16 105
use XNOR2X1  XNOR2X1_37
timestamp 1681708930
transform -1 0 1936 0 1 1170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_38
timestamp 1681708930
transform -1 0 1992 0 1 1170
box -8 -3 64 105
use FILL  FILL_965
timestamp 1681708930
transform 1 0 1992 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_2215
timestamp 1681708930
transform 1 0 2012 0 1 1175
box -3 -3 3 3
use FILL  FILL_966
timestamp 1681708930
transform 1 0 2000 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_50
timestamp 1681708930
transform 1 0 2008 0 1 1170
box -8 -3 46 105
use FILL  FILL_967
timestamp 1681708930
transform 1 0 2048 0 1 1170
box -8 -3 16 105
use FILL  FILL_968
timestamp 1681708930
transform 1 0 2056 0 1 1170
box -8 -3 16 105
use XOR2X1  XOR2X1_113
timestamp 1681708930
transform -1 0 2120 0 1 1170
box -8 -3 64 105
use FILL  FILL_969
timestamp 1681708930
transform 1 0 2120 0 1 1170
box -8 -3 16 105
use FILL  FILL_970
timestamp 1681708930
transform 1 0 2128 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_51
timestamp 1681708930
transform -1 0 2176 0 1 1170
box -8 -3 46 105
use FILL  FILL_971
timestamp 1681708930
transform 1 0 2176 0 1 1170
box -8 -3 16 105
use FILL  FILL_972
timestamp 1681708930
transform 1 0 2184 0 1 1170
box -8 -3 16 105
use FILL  FILL_973
timestamp 1681708930
transform 1 0 2192 0 1 1170
box -8 -3 16 105
use FILL  FILL_974
timestamp 1681708930
transform 1 0 2200 0 1 1170
box -8 -3 16 105
use FILL  FILL_975
timestamp 1681708930
transform 1 0 2208 0 1 1170
box -8 -3 16 105
use FILL  FILL_976
timestamp 1681708930
transform 1 0 2216 0 1 1170
box -8 -3 16 105
use FILL  FILL_977
timestamp 1681708930
transform 1 0 2224 0 1 1170
box -8 -3 16 105
use FILL  FILL_978
timestamp 1681708930
transform 1 0 2232 0 1 1170
box -8 -3 16 105
use FILL  FILL_979
timestamp 1681708930
transform 1 0 2240 0 1 1170
box -8 -3 16 105
use FILL  FILL_980
timestamp 1681708930
transform 1 0 2248 0 1 1170
box -8 -3 16 105
use FILL  FILL_981
timestamp 1681708930
transform 1 0 2256 0 1 1170
box -8 -3 16 105
use FILL  FILL_982
timestamp 1681708930
transform 1 0 2264 0 1 1170
box -8 -3 16 105
use FILL  FILL_983
timestamp 1681708930
transform 1 0 2272 0 1 1170
box -8 -3 16 105
use XOR2X1  XOR2X1_114
timestamp 1681708930
transform 1 0 2280 0 1 1170
box -8 -3 64 105
use FILL  FILL_984
timestamp 1681708930
transform 1 0 2336 0 1 1170
box -8 -3 16 105
use FILL  FILL_985
timestamp 1681708930
transform 1 0 2344 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_159
timestamp 1681708930
transform 1 0 2352 0 1 1170
box -9 -3 26 105
use FILL  FILL_986
timestamp 1681708930
transform 1 0 2368 0 1 1170
box -8 -3 16 105
use FILL  FILL_987
timestamp 1681708930
transform 1 0 2376 0 1 1170
box -8 -3 16 105
use FILL  FILL_988
timestamp 1681708930
transform 1 0 2384 0 1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_61
timestamp 1681708930
transform -1 0 2424 0 1 1170
box -8 -3 34 105
use FILL  FILL_989
timestamp 1681708930
transform 1 0 2424 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_52
timestamp 1681708930
transform -1 0 2472 0 1 1170
box -8 -3 46 105
use INVX2  INVX2_160
timestamp 1681708930
transform -1 0 2488 0 1 1170
box -9 -3 26 105
use FILL  FILL_990
timestamp 1681708930
transform 1 0 2488 0 1 1170
box -8 -3 16 105
use FILL  FILL_1002
timestamp 1681708930
transform 1 0 2496 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_2216
timestamp 1681708930
transform 1 0 2516 0 1 1175
box -3 -3 3 3
use NOR2X1  NOR2X1_54
timestamp 1681708930
transform 1 0 2504 0 1 1170
box -8 -3 32 105
use NAND3X1  NAND3X1_90
timestamp 1681708930
transform 1 0 2528 0 1 1170
box -8 -3 40 105
use FILL  FILL_1003
timestamp 1681708930
transform 1 0 2560 0 1 1170
box -8 -3 16 105
use FILL  FILL_1004
timestamp 1681708930
transform 1 0 2568 0 1 1170
box -8 -3 16 105
use AOI21X1  AOI21X1_34
timestamp 1681708930
transform -1 0 2608 0 1 1170
box -7 -3 39 105
use FILL  FILL_1005
timestamp 1681708930
transform 1 0 2608 0 1 1170
box -8 -3 16 105
use FILL  FILL_1006
timestamp 1681708930
transform 1 0 2616 0 1 1170
box -8 -3 16 105
use FILL  FILL_1007
timestamp 1681708930
transform 1 0 2624 0 1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_55
timestamp 1681708930
transform -1 0 2656 0 1 1170
box -8 -3 32 105
use FILL  FILL_1008
timestamp 1681708930
transform 1 0 2656 0 1 1170
box -8 -3 16 105
use top_mod_new_VIA0  top_mod_new_VIA0_29
timestamp 1681708930
transform 1 0 2688 0 1 1170
box -10 -3 10 3
use M2_M1  M2_M1_2328
timestamp 1681708930
transform 1 0 84 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_2304
timestamp 1681708930
transform 1 0 68 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2305
timestamp 1681708930
transform 1 0 84 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_2385
timestamp 1681708930
transform 1 0 132 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2306
timestamp 1681708930
transform 1 0 164 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2217
timestamp 1681708930
transform 1 0 268 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2218
timestamp 1681708930
transform 1 0 380 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2241
timestamp 1681708930
transform 1 0 284 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2242
timestamp 1681708930
transform 1 0 316 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2243
timestamp 1681708930
transform 1 0 372 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_2329
timestamp 1681708930
transform 1 0 268 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2386
timestamp 1681708930
transform 1 0 172 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2387
timestamp 1681708930
transform 1 0 180 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2388
timestamp 1681708930
transform 1 0 188 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2389
timestamp 1681708930
transform 1 0 244 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2389
timestamp 1681708930
transform 1 0 164 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2390
timestamp 1681708930
transform 1 0 180 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2273
timestamp 1681708930
transform 1 0 340 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_2330
timestamp 1681708930
transform 1 0 292 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2331
timestamp 1681708930
transform 1 0 380 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_2307
timestamp 1681708930
transform 1 0 292 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2274
timestamp 1681708930
transform 1 0 404 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_2332
timestamp 1681708930
transform 1 0 404 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_2294
timestamp 1681708930
transform 1 0 420 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_2390
timestamp 1681708930
transform 1 0 316 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2391
timestamp 1681708930
transform 1 0 372 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2392
timestamp 1681708930
transform 1 0 396 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2362
timestamp 1681708930
transform 1 0 284 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2363
timestamp 1681708930
transform 1 0 324 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2391
timestamp 1681708930
transform 1 0 348 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2392
timestamp 1681708930
transform 1 0 372 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2308
timestamp 1681708930
transform 1 0 412 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2219
timestamp 1681708930
transform 1 0 460 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2244
timestamp 1681708930
transform 1 0 452 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_2321
timestamp 1681708930
transform 1 0 444 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2333
timestamp 1681708930
transform 1 0 436 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_2295
timestamp 1681708930
transform 1 0 444 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_2393
timestamp 1681708930
transform 1 0 420 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2394
timestamp 1681708930
transform 1 0 428 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2364
timestamp 1681708930
transform 1 0 420 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2309
timestamp 1681708930
transform 1 0 444 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2330
timestamp 1681708930
transform 1 0 436 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2275
timestamp 1681708930
transform 1 0 476 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2296
timestamp 1681708930
transform 1 0 468 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_2334
timestamp 1681708930
transform 1 0 476 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2395
timestamp 1681708930
transform 1 0 460 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2396
timestamp 1681708930
transform 1 0 468 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2331
timestamp 1681708930
transform 1 0 460 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2220
timestamp 1681708930
transform 1 0 492 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2245
timestamp 1681708930
transform 1 0 492 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2246
timestamp 1681708930
transform 1 0 524 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2276
timestamp 1681708930
transform 1 0 500 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_2335
timestamp 1681708930
transform 1 0 492 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2336
timestamp 1681708930
transform 1 0 500 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_2297
timestamp 1681708930
transform 1 0 508 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_2322
timestamp 1681708930
transform 1 0 540 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2337
timestamp 1681708930
transform 1 0 524 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2338
timestamp 1681708930
transform 1 0 532 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_2310
timestamp 1681708930
transform 1 0 492 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_2397
timestamp 1681708930
transform 1 0 500 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2398
timestamp 1681708930
transform 1 0 516 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2332
timestamp 1681708930
transform 1 0 500 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2333
timestamp 1681708930
transform 1 0 524 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2365
timestamp 1681708930
transform 1 0 484 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2298
timestamp 1681708930
transform 1 0 540 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_2399
timestamp 1681708930
transform 1 0 540 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2334
timestamp 1681708930
transform 1 0 540 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2299
timestamp 1681708930
transform 1 0 572 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_2400
timestamp 1681708930
transform 1 0 564 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2401
timestamp 1681708930
transform 1 0 572 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2335
timestamp 1681708930
transform 1 0 572 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2376
timestamp 1681708930
transform 1 0 572 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2221
timestamp 1681708930
transform 1 0 596 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2247
timestamp 1681708930
transform 1 0 588 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2277
timestamp 1681708930
transform 1 0 588 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_2339
timestamp 1681708930
transform 1 0 612 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2447
timestamp 1681708930
transform 1 0 612 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_2222
timestamp 1681708930
transform 1 0 644 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2248
timestamp 1681708930
transform 1 0 636 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2300
timestamp 1681708930
transform 1 0 652 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_2340
timestamp 1681708930
transform 1 0 660 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2402
timestamp 1681708930
transform 1 0 636 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2403
timestamp 1681708930
transform 1 0 652 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2336
timestamp 1681708930
transform 1 0 636 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_2448
timestamp 1681708930
transform 1 0 644 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2459
timestamp 1681708930
transform 1 0 628 0 1 1105
box -2 -2 2 2
use M3_M2  M3_M2_2377
timestamp 1681708930
transform 1 0 628 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_2404
timestamp 1681708930
transform 1 0 668 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2337
timestamp 1681708930
transform 1 0 668 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2378
timestamp 1681708930
transform 1 0 660 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2249
timestamp 1681708930
transform 1 0 692 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2250
timestamp 1681708930
transform 1 0 772 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2251
timestamp 1681708930
transform 1 0 788 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2278
timestamp 1681708930
transform 1 0 748 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2279
timestamp 1681708930
transform 1 0 764 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_2341
timestamp 1681708930
transform 1 0 732 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_2301
timestamp 1681708930
transform 1 0 740 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2311
timestamp 1681708930
transform 1 0 732 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_2405
timestamp 1681708930
transform 1 0 740 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2338
timestamp 1681708930
transform 1 0 740 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2223
timestamp 1681708930
transform 1 0 860 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2252
timestamp 1681708930
transform 1 0 852 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_2342
timestamp 1681708930
transform 1 0 756 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2343
timestamp 1681708930
transform 1 0 764 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2344
timestamp 1681708930
transform 1 0 812 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2345
timestamp 1681708930
transform 1 0 820 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_2312
timestamp 1681708930
transform 1 0 756 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_2406
timestamp 1681708930
transform 1 0 764 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2313
timestamp 1681708930
transform 1 0 788 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2314
timestamp 1681708930
transform 1 0 820 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_2407
timestamp 1681708930
transform 1 0 844 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2366
timestamp 1681708930
transform 1 0 748 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2379
timestamp 1681708930
transform 1 0 732 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2224
timestamp 1681708930
transform 1 0 892 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2280
timestamp 1681708930
transform 1 0 884 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_2346
timestamp 1681708930
transform 1 0 884 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2408
timestamp 1681708930
transform 1 0 876 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2339
timestamp 1681708930
transform 1 0 836 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2340
timestamp 1681708930
transform 1 0 868 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2367
timestamp 1681708930
transform 1 0 844 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2380
timestamp 1681708930
transform 1 0 812 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2381
timestamp 1681708930
transform 1 0 844 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2281
timestamp 1681708930
transform 1 0 940 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_2409
timestamp 1681708930
transform 1 0 916 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2410
timestamp 1681708930
transform 1 0 940 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2341
timestamp 1681708930
transform 1 0 892 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2342
timestamp 1681708930
transform 1 0 916 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2253
timestamp 1681708930
transform 1 0 972 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_2347
timestamp 1681708930
transform 1 0 964 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2348
timestamp 1681708930
transform 1 0 972 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_2315
timestamp 1681708930
transform 1 0 964 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2225
timestamp 1681708930
transform 1 0 1012 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2226
timestamp 1681708930
transform 1 0 1036 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_2319
timestamp 1681708930
transform 1 0 1036 0 1 1155
box -2 -2 2 2
use M2_M1  M2_M1_2323
timestamp 1681708930
transform 1 0 1036 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_2227
timestamp 1681708930
transform 1 0 1060 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_2320
timestamp 1681708930
transform 1 0 1060 0 1 1155
box -2 -2 2 2
use M2_M1  M2_M1_2324
timestamp 1681708930
transform 1 0 1052 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2349
timestamp 1681708930
transform 1 0 1052 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_2316
timestamp 1681708930
transform 1 0 1060 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_2350
timestamp 1681708930
transform 1 0 1076 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2351
timestamp 1681708930
transform 1 0 1092 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2411
timestamp 1681708930
transform 1 0 1084 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2412
timestamp 1681708930
transform 1 0 1100 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2343
timestamp 1681708930
transform 1 0 1084 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2368
timestamp 1681708930
transform 1 0 1076 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_2413
timestamp 1681708930
transform 1 0 1116 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2352
timestamp 1681708930
transform 1 0 1124 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_2344
timestamp 1681708930
transform 1 0 1116 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2228
timestamp 1681708930
transform 1 0 1140 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_2353
timestamp 1681708930
transform 1 0 1164 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2354
timestamp 1681708930
transform 1 0 1212 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2414
timestamp 1681708930
transform 1 0 1204 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2449
timestamp 1681708930
transform 1 0 1212 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_2369
timestamp 1681708930
transform 1 0 1212 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2282
timestamp 1681708930
transform 1 0 1260 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2317
timestamp 1681708930
transform 1 0 1308 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2370
timestamp 1681708930
transform 1 0 1308 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2393
timestamp 1681708930
transform 1 0 1300 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2229
timestamp 1681708930
transform 1 0 1348 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2254
timestamp 1681708930
transform 1 0 1380 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_2415
timestamp 1681708930
transform 1 0 1372 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2255
timestamp 1681708930
transform 1 0 1396 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_2355
timestamp 1681708930
transform 1 0 1388 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_2382
timestamp 1681708930
transform 1 0 1388 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2394
timestamp 1681708930
transform 1 0 1396 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2302
timestamp 1681708930
transform 1 0 1460 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_2416
timestamp 1681708930
transform 1 0 1492 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2345
timestamp 1681708930
transform 1 0 1492 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2256
timestamp 1681708930
transform 1 0 1508 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_2450
timestamp 1681708930
transform 1 0 1500 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2451
timestamp 1681708930
transform 1 0 1508 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2460
timestamp 1681708930
transform 1 0 1524 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_2356
timestamp 1681708930
transform 1 0 1564 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2417
timestamp 1681708930
transform 1 0 1548 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2318
timestamp 1681708930
transform 1 0 1564 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2346
timestamp 1681708930
transform 1 0 1548 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_2452
timestamp 1681708930
transform 1 0 1556 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2461
timestamp 1681708930
transform 1 0 1540 0 1 1105
box -2 -2 2 2
use M3_M2  M3_M2_2257
timestamp 1681708930
transform 1 0 1612 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2258
timestamp 1681708930
transform 1 0 1636 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2259
timestamp 1681708930
transform 1 0 1652 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_2357
timestamp 1681708930
transform 1 0 1612 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2358
timestamp 1681708930
transform 1 0 1620 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_2230
timestamp 1681708930
transform 1 0 1732 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2283
timestamp 1681708930
transform 1 0 1684 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2284
timestamp 1681708930
transform 1 0 1716 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2285
timestamp 1681708930
transform 1 0 1732 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_2359
timestamp 1681708930
transform 1 0 1668 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2360
timestamp 1681708930
transform 1 0 1684 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_2260
timestamp 1681708930
transform 1 0 1780 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_2418
timestamp 1681708930
transform 1 0 1620 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2419
timestamp 1681708930
transform 1 0 1644 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2319
timestamp 1681708930
transform 1 0 1668 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_2420
timestamp 1681708930
transform 1 0 1732 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2320
timestamp 1681708930
transform 1 0 1756 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_2421
timestamp 1681708930
transform 1 0 1764 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2422
timestamp 1681708930
transform 1 0 1772 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2347
timestamp 1681708930
transform 1 0 1732 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2348
timestamp 1681708930
transform 1 0 1772 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2395
timestamp 1681708930
transform 1 0 1676 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2396
timestamp 1681708930
transform 1 0 1708 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2261
timestamp 1681708930
transform 1 0 1796 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_2423
timestamp 1681708930
transform 1 0 1796 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2349
timestamp 1681708930
transform 1 0 1796 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2262
timestamp 1681708930
transform 1 0 1836 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2231
timestamp 1681708930
transform 1 0 1868 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2263
timestamp 1681708930
transform 1 0 1884 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_2361
timestamp 1681708930
transform 1 0 1812 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2362
timestamp 1681708930
transform 1 0 1820 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2363
timestamp 1681708930
transform 1 0 1836 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2364
timestamp 1681708930
transform 1 0 1844 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2424
timestamp 1681708930
transform 1 0 1828 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2321
timestamp 1681708930
transform 1 0 1844 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2232
timestamp 1681708930
transform 1 0 1908 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_2365
timestamp 1681708930
transform 1 0 1900 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2425
timestamp 1681708930
transform 1 0 1852 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2426
timestamp 1681708930
transform 1 0 1876 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2350
timestamp 1681708930
transform 1 0 1852 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2351
timestamp 1681708930
transform 1 0 1876 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2286
timestamp 1681708930
transform 1 0 1916 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_2366
timestamp 1681708930
transform 1 0 1916 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_2233
timestamp 1681708930
transform 1 0 2028 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2264
timestamp 1681708930
transform 1 0 1972 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2265
timestamp 1681708930
transform 1 0 1988 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2266
timestamp 1681708930
transform 1 0 2004 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_2367
timestamp 1681708930
transform 1 0 1964 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2368
timestamp 1681708930
transform 1 0 1972 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2427
timestamp 1681708930
transform 1 0 1940 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2234
timestamp 1681708930
transform 1 0 2084 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2235
timestamp 1681708930
transform 1 0 2116 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2236
timestamp 1681708930
transform 1 0 2140 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2267
timestamp 1681708930
transform 1 0 2068 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_2369
timestamp 1681708930
transform 1 0 2020 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2370
timestamp 1681708930
transform 1 0 2028 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2428
timestamp 1681708930
transform 1 0 1988 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2322
timestamp 1681708930
transform 1 0 1996 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_2429
timestamp 1681708930
transform 1 0 2020 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2352
timestamp 1681708930
transform 1 0 1964 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2371
timestamp 1681708930
transform 1 0 1924 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2383
timestamp 1681708930
transform 1 0 1932 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2397
timestamp 1681708930
transform 1 0 1916 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2353
timestamp 1681708930
transform 1 0 2020 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2372
timestamp 1681708930
transform 1 0 2012 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2268
timestamp 1681708930
transform 1 0 2124 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_2371
timestamp 1681708930
transform 1 0 2076 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2372
timestamp 1681708930
transform 1 0 2084 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_2287
timestamp 1681708930
transform 1 0 2156 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2288
timestamp 1681708930
transform 1 0 2172 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_2373
timestamp 1681708930
transform 1 0 2132 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2374
timestamp 1681708930
transform 1 0 2140 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2375
timestamp 1681708930
transform 1 0 2148 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2376
timestamp 1681708930
transform 1 0 2164 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2377
timestamp 1681708930
transform 1 0 2172 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_2323
timestamp 1681708930
transform 1 0 2084 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2324
timestamp 1681708930
transform 1 0 2100 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_2430
timestamp 1681708930
transform 1 0 2108 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2237
timestamp 1681708930
transform 1 0 2284 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2289
timestamp 1681708930
transform 1 0 2276 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_2378
timestamp 1681708930
transform 1 0 2204 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2431
timestamp 1681708930
transform 1 0 2156 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2432
timestamp 1681708930
transform 1 0 2172 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2433
timestamp 1681708930
transform 1 0 2188 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2434
timestamp 1681708930
transform 1 0 2228 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2325
timestamp 1681708930
transform 1 0 2268 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2269
timestamp 1681708930
transform 1 0 2348 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_2379
timestamp 1681708930
transform 1 0 2340 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2435
timestamp 1681708930
transform 1 0 2284 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2354
timestamp 1681708930
transform 1 0 2188 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2355
timestamp 1681708930
transform 1 0 2228 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2384
timestamp 1681708930
transform 1 0 2276 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2326
timestamp 1681708930
transform 1 0 2308 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_2436
timestamp 1681708930
transform 1 0 2316 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2437
timestamp 1681708930
transform 1 0 2372 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2453
timestamp 1681708930
transform 1 0 2356 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_2373
timestamp 1681708930
transform 1 0 2348 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2356
timestamp 1681708930
transform 1 0 2372 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_2454
timestamp 1681708930
transform 1 0 2380 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2462
timestamp 1681708930
transform 1 0 2372 0 1 1105
box -2 -2 2 2
use M3_M2  M3_M2_2374
timestamp 1681708930
transform 1 0 2380 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2270
timestamp 1681708930
transform 1 0 2404 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2290
timestamp 1681708930
transform 1 0 2404 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2238
timestamp 1681708930
transform 1 0 2428 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_2380
timestamp 1681708930
transform 1 0 2404 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_2327
timestamp 1681708930
transform 1 0 2396 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_2467
timestamp 1681708930
transform 1 0 2388 0 1 1095
box -2 -2 2 2
use M3_M2  M3_M2_2398
timestamp 1681708930
transform 1 0 2388 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2303
timestamp 1681708930
transform 1 0 2420 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_2463
timestamp 1681708930
transform 1 0 2412 0 1 1105
box -2 -2 2 2
use M3_M2  M3_M2_2385
timestamp 1681708930
transform 1 0 2412 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_2438
timestamp 1681708930
transform 1 0 2428 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2291
timestamp 1681708930
transform 1 0 2436 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2328
timestamp 1681708930
transform 1 0 2436 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2357
timestamp 1681708930
transform 1 0 2428 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_2455
timestamp 1681708930
transform 1 0 2436 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_2239
timestamp 1681708930
transform 1 0 2452 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_2325
timestamp 1681708930
transform 1 0 2460 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_2399
timestamp 1681708930
transform 1 0 2452 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2271
timestamp 1681708930
transform 1 0 2484 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2292
timestamp 1681708930
transform 1 0 2476 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_2381
timestamp 1681708930
transform 1 0 2484 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2439
timestamp 1681708930
transform 1 0 2476 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2386
timestamp 1681708930
transform 1 0 2476 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2400
timestamp 1681708930
transform 1 0 2476 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_2382
timestamp 1681708930
transform 1 0 2500 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_2329
timestamp 1681708930
transform 1 0 2500 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_2440
timestamp 1681708930
transform 1 0 2508 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2441
timestamp 1681708930
transform 1 0 2516 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2240
timestamp 1681708930
transform 1 0 2532 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2272
timestamp 1681708930
transform 1 0 2572 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_2326
timestamp 1681708930
transform 1 0 2572 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2383
timestamp 1681708930
transform 1 0 2588 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2442
timestamp 1681708930
transform 1 0 2556 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2443
timestamp 1681708930
transform 1 0 2572 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2358
timestamp 1681708930
transform 1 0 2556 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_2456
timestamp 1681708930
transform 1 0 2564 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2464
timestamp 1681708930
transform 1 0 2548 0 1 1105
box -2 -2 2 2
use M3_M2  M3_M2_2293
timestamp 1681708930
transform 1 0 2628 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_2327
timestamp 1681708930
transform 1 0 2636 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2384
timestamp 1681708930
transform 1 0 2636 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2444
timestamp 1681708930
transform 1 0 2596 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2445
timestamp 1681708930
transform 1 0 2620 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2359
timestamp 1681708930
transform 1 0 2596 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_2457
timestamp 1681708930
transform 1 0 2604 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_2360
timestamp 1681708930
transform 1 0 2620 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_2458
timestamp 1681708930
transform 1 0 2628 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_2361
timestamp 1681708930
transform 1 0 2636 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2375
timestamp 1681708930
transform 1 0 2604 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_2465
timestamp 1681708930
transform 1 0 2612 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_2466
timestamp 1681708930
transform 1 0 2620 0 1 1105
box -2 -2 2 2
use M3_M2  M3_M2_2387
timestamp 1681708930
transform 1 0 2612 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2401
timestamp 1681708930
transform 1 0 2620 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_2446
timestamp 1681708930
transform 1 0 2652 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_2388
timestamp 1681708930
transform 1 0 2644 0 1 1095
box -3 -3 3 3
use top_mod_new_VIA0  top_mod_new_VIA0_30
timestamp 1681708930
transform 1 0 24 0 1 1070
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_59
timestamp 1681708930
transform 1 0 72 0 -1 1170
box -8 -3 104 105
use INVX2  INVX2_152
timestamp 1681708930
transform 1 0 168 0 -1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_60
timestamp 1681708930
transform -1 0 280 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_61
timestamp 1681708930
transform 1 0 280 0 -1 1170
box -8 -3 104 105
use BUFX2  BUFX2_4
timestamp 1681708930
transform -1 0 400 0 -1 1170
box -5 -3 28 105
use BUFX2  BUFX2_5
timestamp 1681708930
transform -1 0 424 0 -1 1170
box -5 -3 28 105
use INVX2  INVX2_153
timestamp 1681708930
transform -1 0 440 0 -1 1170
box -9 -3 26 105
use NOR2X1  NOR2X1_51
timestamp 1681708930
transform 1 0 440 0 -1 1170
box -8 -3 32 105
use FILL  FILL_892
timestamp 1681708930
transform 1 0 464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_893
timestamp 1681708930
transform 1 0 472 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_154
timestamp 1681708930
transform -1 0 496 0 -1 1170
box -9 -3 26 105
use AOI22X1  AOI22X1_48
timestamp 1681708930
transform 1 0 496 0 -1 1170
box -8 -3 46 105
use FILL  FILL_894
timestamp 1681708930
transform 1 0 536 0 -1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_52
timestamp 1681708930
transform 1 0 544 0 -1 1170
box -8 -3 32 105
use FILL  FILL_895
timestamp 1681708930
transform 1 0 568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_896
timestamp 1681708930
transform 1 0 576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_897
timestamp 1681708930
transform 1 0 584 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_155
timestamp 1681708930
transform -1 0 608 0 -1 1170
box -9 -3 26 105
use FILL  FILL_898
timestamp 1681708930
transform 1 0 608 0 -1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_84
timestamp 1681708930
transform -1 0 648 0 -1 1170
box -8 -3 40 105
use M3_M2  M3_M2_2402
timestamp 1681708930
transform 1 0 668 0 1 1075
box -3 -3 3 3
use INVX2  INVX2_156
timestamp 1681708930
transform -1 0 664 0 -1 1170
box -9 -3 26 105
use FILL  FILL_899
timestamp 1681708930
transform 1 0 664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_900
timestamp 1681708930
transform 1 0 672 0 -1 1170
box -8 -3 16 105
use XNOR2X1  XNOR2X1_36
timestamp 1681708930
transform -1 0 736 0 -1 1170
box -8 -3 64 105
use M3_M2  M3_M2_2403
timestamp 1681708930
transform 1 0 748 0 1 1075
box -3 -3 3 3
use BUFX2  BUFX2_6
timestamp 1681708930
transform 1 0 736 0 -1 1170
box -5 -3 28 105
use XOR2X1  XOR2X1_107
timestamp 1681708930
transform -1 0 816 0 -1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_108
timestamp 1681708930
transform 1 0 816 0 -1 1170
box -8 -3 64 105
use FILL  FILL_901
timestamp 1681708930
transform 1 0 872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_902
timestamp 1681708930
transform 1 0 880 0 -1 1170
box -8 -3 16 105
use XOR2X1  XOR2X1_109
timestamp 1681708930
transform 1 0 888 0 -1 1170
box -8 -3 64 105
use FILL  FILL_903
timestamp 1681708930
transform 1 0 944 0 -1 1170
box -8 -3 16 105
use FILL  FILL_904
timestamp 1681708930
transform 1 0 952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_905
timestamp 1681708930
transform 1 0 960 0 -1 1170
box -8 -3 16 105
use FILL  FILL_906
timestamp 1681708930
transform 1 0 968 0 -1 1170
box -8 -3 16 105
use XOR2X1  XOR2X1_110
timestamp 1681708930
transform -1 0 1032 0 -1 1170
box -8 -3 64 105
use FILL  FILL_907
timestamp 1681708930
transform 1 0 1032 0 -1 1170
box -8 -3 16 105
use FILL  FILL_908
timestamp 1681708930
transform 1 0 1040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_909
timestamp 1681708930
transform 1 0 1048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_910
timestamp 1681708930
transform 1 0 1056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_911
timestamp 1681708930
transform 1 0 1064 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_22
timestamp 1681708930
transform 1 0 1072 0 -1 1170
box -8 -3 46 105
use FILL  FILL_912
timestamp 1681708930
transform 1 0 1112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_913
timestamp 1681708930
transform 1 0 1120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_914
timestamp 1681708930
transform 1 0 1128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_915
timestamp 1681708930
transform 1 0 1136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_916
timestamp 1681708930
transform 1 0 1144 0 -1 1170
box -8 -3 16 105
use FILL  FILL_917
timestamp 1681708930
transform 1 0 1152 0 -1 1170
box -8 -3 16 105
use FILL  FILL_918
timestamp 1681708930
transform 1 0 1160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_919
timestamp 1681708930
transform 1 0 1168 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_157
timestamp 1681708930
transform 1 0 1176 0 -1 1170
box -9 -3 26 105
use NAND2X1  NAND2X1_58
timestamp 1681708930
transform 1 0 1192 0 -1 1170
box -8 -3 32 105
use FILL  FILL_920
timestamp 1681708930
transform 1 0 1216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_921
timestamp 1681708930
transform 1 0 1224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_922
timestamp 1681708930
transform 1 0 1232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_923
timestamp 1681708930
transform 1 0 1240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_924
timestamp 1681708930
transform 1 0 1248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_925
timestamp 1681708930
transform 1 0 1256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_926
timestamp 1681708930
transform 1 0 1264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_927
timestamp 1681708930
transform 1 0 1272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_928
timestamp 1681708930
transform 1 0 1280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_929
timestamp 1681708930
transform 1 0 1288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_930
timestamp 1681708930
transform 1 0 1296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_931
timestamp 1681708930
transform 1 0 1304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_932
timestamp 1681708930
transform 1 0 1312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_933
timestamp 1681708930
transform 1 0 1320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_934
timestamp 1681708930
transform 1 0 1328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_935
timestamp 1681708930
transform 1 0 1336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_936
timestamp 1681708930
transform 1 0 1344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_937
timestamp 1681708930
transform 1 0 1352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_938
timestamp 1681708930
transform 1 0 1360 0 -1 1170
box -8 -3 16 105
use FILL  FILL_939
timestamp 1681708930
transform 1 0 1368 0 -1 1170
box -8 -3 16 105
use FILL  FILL_940
timestamp 1681708930
transform 1 0 1376 0 -1 1170
box -8 -3 16 105
use XOR2X1  XOR2X1_111
timestamp 1681708930
transform -1 0 1440 0 -1 1170
box -8 -3 64 105
use FILL  FILL_941
timestamp 1681708930
transform 1 0 1440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_942
timestamp 1681708930
transform 1 0 1448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_943
timestamp 1681708930
transform 1 0 1456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_946
timestamp 1681708930
transform 1 0 1464 0 -1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_86
timestamp 1681708930
transform -1 0 1504 0 -1 1170
box -8 -3 40 105
use FILL  FILL_947
timestamp 1681708930
transform 1 0 1504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_949
timestamp 1681708930
transform 1 0 1512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_991
timestamp 1681708930
transform 1 0 1520 0 -1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_87
timestamp 1681708930
transform -1 0 1560 0 -1 1170
box -8 -3 40 105
use XOR2X1  XOR2X1_115
timestamp 1681708930
transform 1 0 1560 0 -1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_116
timestamp 1681708930
transform 1 0 1616 0 -1 1170
box -8 -3 64 105
use DFFNEGX1  DFFNEGX1_63
timestamp 1681708930
transform 1 0 1672 0 -1 1170
box -8 -3 104 105
use INVX2  INVX2_161
timestamp 1681708930
transform -1 0 1784 0 -1 1170
box -9 -3 26 105
use FILL  FILL_992
timestamp 1681708930
transform 1 0 1784 0 -1 1170
box -8 -3 16 105
use FILL  FILL_993
timestamp 1681708930
transform 1 0 1792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_994
timestamp 1681708930
transform 1 0 1800 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_2404
timestamp 1681708930
transform 1 0 1844 0 1 1075
box -3 -3 3 3
use AOI22X1  AOI22X1_53
timestamp 1681708930
transform -1 0 1848 0 -1 1170
box -8 -3 46 105
use XOR2X1  XOR2X1_117
timestamp 1681708930
transform 1 0 1848 0 -1 1170
box -8 -3 64 105
use FILL  FILL_995
timestamp 1681708930
transform 1 0 1904 0 -1 1170
box -8 -3 16 105
use XOR2X1  XOR2X1_118
timestamp 1681708930
transform 1 0 1912 0 -1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_119
timestamp 1681708930
transform -1 0 2024 0 -1 1170
box -8 -3 64 105
use M3_M2  M3_M2_2405
timestamp 1681708930
transform 1 0 2100 0 1 1075
box -3 -3 3 3
use XNOR2X1  XNOR2X1_39
timestamp 1681708930
transform -1 0 2080 0 -1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_120
timestamp 1681708930
transform -1 0 2136 0 -1 1170
box -8 -3 64 105
use M3_M2  M3_M2_2406
timestamp 1681708930
transform 1 0 2164 0 1 1075
box -3 -3 3 3
use AOI22X1  AOI22X1_54
timestamp 1681708930
transform -1 0 2176 0 -1 1170
box -8 -3 46 105
use M3_M2  M3_M2_2407
timestamp 1681708930
transform 1 0 2204 0 1 1075
box -3 -3 3 3
use INVX2  INVX2_162
timestamp 1681708930
transform 1 0 2176 0 -1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_64
timestamp 1681708930
transform 1 0 2192 0 -1 1170
box -8 -3 104 105
use XOR2X1  XOR2X1_121
timestamp 1681708930
transform -1 0 2344 0 -1 1170
box -8 -3 64 105
use FILL  FILL_996
timestamp 1681708930
transform 1 0 2344 0 -1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_88
timestamp 1681708930
transform -1 0 2384 0 -1 1170
box -8 -3 40 105
use FILL  FILL_997
timestamp 1681708930
transform 1 0 2384 0 -1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_89
timestamp 1681708930
transform 1 0 2392 0 -1 1170
box -8 -3 40 105
use FILL  FILL_998
timestamp 1681708930
transform 1 0 2424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_999
timestamp 1681708930
transform 1 0 2432 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_163
timestamp 1681708930
transform -1 0 2456 0 -1 1170
box -9 -3 26 105
use NOR2X1  NOR2X1_53
timestamp 1681708930
transform 1 0 2456 0 -1 1170
box -8 -3 32 105
use FILL  FILL_1000
timestamp 1681708930
transform 1 0 2480 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1001
timestamp 1681708930
transform 1 0 2488 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_164
timestamp 1681708930
transform 1 0 2496 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_165
timestamp 1681708930
transform -1 0 2528 0 -1 1170
box -9 -3 26 105
use FILL  FILL_1009
timestamp 1681708930
transform 1 0 2528 0 -1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_91
timestamp 1681708930
transform -1 0 2568 0 -1 1170
box -8 -3 40 105
use AOI21X1  AOI21X1_35
timestamp 1681708930
transform -1 0 2600 0 -1 1170
box -7 -3 39 105
use NAND3X1  NAND3X1_92
timestamp 1681708930
transform -1 0 2632 0 -1 1170
box -8 -3 40 105
use NOR2X1  NOR2X1_56
timestamp 1681708930
transform 1 0 2632 0 -1 1170
box -8 -3 32 105
use FILL  FILL_1010
timestamp 1681708930
transform 1 0 2656 0 -1 1170
box -8 -3 16 105
use top_mod_new_VIA0  top_mod_new_VIA0_31
timestamp 1681708930
transform 1 0 2712 0 1 1070
box -10 -3 10 3
use M3_M2  M3_M2_2467
timestamp 1681708930
transform 1 0 132 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2483
timestamp 1681708930
transform 1 0 68 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_2501
timestamp 1681708930
transform 1 0 76 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2502
timestamp 1681708930
transform 1 0 108 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2424
timestamp 1681708930
transform 1 0 164 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_2471
timestamp 1681708930
transform 1 0 148 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_2468
timestamp 1681708930
transform 1 0 156 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2469
timestamp 1681708930
transform 1 0 188 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2484
timestamp 1681708930
transform 1 0 132 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2485
timestamp 1681708930
transform 1 0 140 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2486
timestamp 1681708930
transform 1 0 148 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2487
timestamp 1681708930
transform 1 0 172 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2488
timestamp 1681708930
transform 1 0 188 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2550
timestamp 1681708930
transform 1 0 68 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2551
timestamp 1681708930
transform 1 0 124 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2552
timestamp 1681708930
transform 1 0 132 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2544
timestamp 1681708930
transform 1 0 68 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2545
timestamp 1681708930
transform 1 0 132 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_2638
timestamp 1681708930
transform 1 0 68 0 1 985
box -2 -2 2 2
use M3_M2  M3_M2_2565
timestamp 1681708930
transform 1 0 76 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2566
timestamp 1681708930
transform 1 0 108 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_2553
timestamp 1681708930
transform 1 0 164 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2530
timestamp 1681708930
transform 1 0 172 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_2554
timestamp 1681708930
transform 1 0 180 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2546
timestamp 1681708930
transform 1 0 148 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_2489
timestamp 1681708930
transform 1 0 204 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_2531
timestamp 1681708930
transform 1 0 212 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2425
timestamp 1681708930
transform 1 0 260 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2426
timestamp 1681708930
transform 1 0 292 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2437
timestamp 1681708930
transform 1 0 244 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2438
timestamp 1681708930
transform 1 0 276 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_2468
timestamp 1681708930
transform 1 0 284 0 1 1035
box -2 -2 2 2
use M3_M2  M3_M2_2503
timestamp 1681708930
transform 1 0 236 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_2472
timestamp 1681708930
transform 1 0 276 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2490
timestamp 1681708930
transform 1 0 244 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2491
timestamp 1681708930
transform 1 0 260 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2555
timestamp 1681708930
transform 1 0 220 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2556
timestamp 1681708930
transform 1 0 228 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2557
timestamp 1681708930
transform 1 0 236 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2547
timestamp 1681708930
transform 1 0 204 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_2630
timestamp 1681708930
transform 1 0 212 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_2532
timestamp 1681708930
transform 1 0 244 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2470
timestamp 1681708930
transform 1 0 300 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2473
timestamp 1681708930
transform 1 0 308 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_2504
timestamp 1681708930
transform 1 0 284 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_2492
timestamp 1681708930
transform 1 0 292 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_2505
timestamp 1681708930
transform 1 0 308 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_2474
timestamp 1681708930
transform 1 0 324 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2493
timestamp 1681708930
transform 1 0 316 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2558
timestamp 1681708930
transform 1 0 252 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2559
timestamp 1681708930
transform 1 0 268 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2506
timestamp 1681708930
transform 1 0 324 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_2560
timestamp 1681708930
transform 1 0 308 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2533
timestamp 1681708930
transform 1 0 316 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2548
timestamp 1681708930
transform 1 0 316 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_2561
timestamp 1681708930
transform 1 0 348 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2471
timestamp 1681708930
transform 1 0 356 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2494
timestamp 1681708930
transform 1 0 356 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_2439
timestamp 1681708930
transform 1 0 436 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2472
timestamp 1681708930
transform 1 0 372 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2473
timestamp 1681708930
transform 1 0 404 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2495
timestamp 1681708930
transform 1 0 380 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2496
timestamp 1681708930
transform 1 0 404 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2497
timestamp 1681708930
transform 1 0 428 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2562
timestamp 1681708930
transform 1 0 380 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2549
timestamp 1681708930
transform 1 0 380 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2507
timestamp 1681708930
transform 1 0 452 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_2498
timestamp 1681708930
transform 1 0 460 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2563
timestamp 1681708930
transform 1 0 428 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2564
timestamp 1681708930
transform 1 0 436 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2565
timestamp 1681708930
transform 1 0 452 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2567
timestamp 1681708930
transform 1 0 396 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2534
timestamp 1681708930
transform 1 0 460 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2440
timestamp 1681708930
transform 1 0 508 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2474
timestamp 1681708930
transform 1 0 500 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2499
timestamp 1681708930
transform 1 0 492 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2500
timestamp 1681708930
transform 1 0 500 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2501
timestamp 1681708930
transform 1 0 524 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2566
timestamp 1681708930
transform 1 0 468 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2550
timestamp 1681708930
transform 1 0 452 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2551
timestamp 1681708930
transform 1 0 476 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2568
timestamp 1681708930
transform 1 0 444 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2569
timestamp 1681708930
transform 1 0 468 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_2567
timestamp 1681708930
transform 1 0 532 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2552
timestamp 1681708930
transform 1 0 532 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2408
timestamp 1681708930
transform 1 0 556 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2441
timestamp 1681708930
transform 1 0 564 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_2502
timestamp 1681708930
transform 1 0 564 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2568
timestamp 1681708930
transform 1 0 556 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2569
timestamp 1681708930
transform 1 0 564 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2631
timestamp 1681708930
transform 1 0 540 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_2570
timestamp 1681708930
transform 1 0 524 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2553
timestamp 1681708930
transform 1 0 564 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2427
timestamp 1681708930
transform 1 0 580 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_2475
timestamp 1681708930
transform 1 0 580 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_2475
timestamp 1681708930
transform 1 0 588 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2503
timestamp 1681708930
transform 1 0 596 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_2508
timestamp 1681708930
transform 1 0 604 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2428
timestamp 1681708930
transform 1 0 628 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_2570
timestamp 1681708930
transform 1 0 604 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2571
timestamp 1681708930
transform 1 0 620 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2554
timestamp 1681708930
transform 1 0 620 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2442
timestamp 1681708930
transform 1 0 636 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_2632
timestamp 1681708930
transform 1 0 628 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_2509
timestamp 1681708930
transform 1 0 644 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2476
timestamp 1681708930
transform 1 0 676 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2476
timestamp 1681708930
transform 1 0 700 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2504
timestamp 1681708930
transform 1 0 652 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2505
timestamp 1681708930
transform 1 0 676 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2506
timestamp 1681708930
transform 1 0 692 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_2535
timestamp 1681708930
transform 1 0 652 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_2572
timestamp 1681708930
transform 1 0 660 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2573
timestamp 1681708930
transform 1 0 668 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2536
timestamp 1681708930
transform 1 0 684 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2429
timestamp 1681708930
transform 1 0 716 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_2574
timestamp 1681708930
transform 1 0 708 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2571
timestamp 1681708930
transform 1 0 708 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2409
timestamp 1681708930
transform 1 0 756 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2477
timestamp 1681708930
transform 1 0 732 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2430
timestamp 1681708930
transform 1 0 788 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2431
timestamp 1681708930
transform 1 0 804 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2443
timestamp 1681708930
transform 1 0 780 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2510
timestamp 1681708930
transform 1 0 756 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_2507
timestamp 1681708930
transform 1 0 788 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2575
timestamp 1681708930
transform 1 0 724 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2576
timestamp 1681708930
transform 1 0 732 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2555
timestamp 1681708930
transform 1 0 724 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2511
timestamp 1681708930
transform 1 0 804 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2512
timestamp 1681708930
transform 1 0 820 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_2577
timestamp 1681708930
transform 1 0 780 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2578
timestamp 1681708930
transform 1 0 788 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2556
timestamp 1681708930
transform 1 0 780 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2572
timestamp 1681708930
transform 1 0 764 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2432
timestamp 1681708930
transform 1 0 948 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2444
timestamp 1681708930
transform 1 0 876 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2445
timestamp 1681708930
transform 1 0 900 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2478
timestamp 1681708930
transform 1 0 868 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2508
timestamp 1681708930
transform 1 0 868 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2509
timestamp 1681708930
transform 1 0 876 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2579
timestamp 1681708930
transform 1 0 836 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2580
timestamp 1681708930
transform 1 0 844 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2557
timestamp 1681708930
transform 1 0 844 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2573
timestamp 1681708930
transform 1 0 804 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2513
timestamp 1681708930
transform 1 0 892 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_2510
timestamp 1681708930
transform 1 0 948 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2581
timestamp 1681708930
transform 1 0 892 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2582
timestamp 1681708930
transform 1 0 900 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2583
timestamp 1681708930
transform 1 0 948 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2574
timestamp 1681708930
transform 1 0 900 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2433
timestamp 1681708930
transform 1 0 1028 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2479
timestamp 1681708930
transform 1 0 1004 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2511
timestamp 1681708930
transform 1 0 1004 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2584
timestamp 1681708930
transform 1 0 972 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2585
timestamp 1681708930
transform 1 0 980 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2586
timestamp 1681708930
transform 1 0 1028 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2587
timestamp 1681708930
transform 1 0 1052 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2558
timestamp 1681708930
transform 1 0 1044 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2446
timestamp 1681708930
transform 1 0 1068 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_2477
timestamp 1681708930
transform 1 0 1060 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_2514
timestamp 1681708930
transform 1 0 1060 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_2512
timestamp 1681708930
transform 1 0 1076 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2513
timestamp 1681708930
transform 1 0 1100 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2588
timestamp 1681708930
transform 1 0 1116 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2537
timestamp 1681708930
transform 1 0 1124 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_2633
timestamp 1681708930
transform 1 0 1132 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2589
timestamp 1681708930
transform 1 0 1148 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2480
timestamp 1681708930
transform 1 0 1164 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2514
timestamp 1681708930
transform 1 0 1164 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_2575
timestamp 1681708930
transform 1 0 1180 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_2515
timestamp 1681708930
transform 1 0 1204 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2590
timestamp 1681708930
transform 1 0 1196 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2447
timestamp 1681708930
transform 1 0 1244 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2481
timestamp 1681708930
transform 1 0 1236 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2410
timestamp 1681708930
transform 1 0 1276 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2482
timestamp 1681708930
transform 1 0 1268 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2515
timestamp 1681708930
transform 1 0 1252 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2411
timestamp 1681708930
transform 1 0 1324 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2416
timestamp 1681708930
transform 1 0 1316 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2417
timestamp 1681708930
transform 1 0 1340 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2448
timestamp 1681708930
transform 1 0 1292 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2449
timestamp 1681708930
transform 1 0 1308 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2450
timestamp 1681708930
transform 1 0 1324 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2483
timestamp 1681708930
transform 1 0 1300 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2516
timestamp 1681708930
transform 1 0 1260 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2517
timestamp 1681708930
transform 1 0 1284 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2591
timestamp 1681708930
transform 1 0 1252 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2592
timestamp 1681708930
transform 1 0 1268 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2538
timestamp 1681708930
transform 1 0 1284 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_2518
timestamp 1681708930
transform 1 0 1308 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2593
timestamp 1681708930
transform 1 0 1300 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2594
timestamp 1681708930
transform 1 0 1308 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2634
timestamp 1681708930
transform 1 0 1284 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_2539
timestamp 1681708930
transform 1 0 1316 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_2635
timestamp 1681708930
transform 1 0 1316 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_2576
timestamp 1681708930
transform 1 0 1300 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2451
timestamp 1681708930
transform 1 0 1356 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2452
timestamp 1681708930
transform 1 0 1388 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2484
timestamp 1681708930
transform 1 0 1332 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2519
timestamp 1681708930
transform 1 0 1332 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2520
timestamp 1681708930
transform 1 0 1356 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_2516
timestamp 1681708930
transform 1 0 1372 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_2595
timestamp 1681708930
transform 1 0 1332 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2596
timestamp 1681708930
transform 1 0 1388 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2597
timestamp 1681708930
transform 1 0 1396 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2453
timestamp 1681708930
transform 1 0 1484 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2454
timestamp 1681708930
transform 1 0 1500 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2485
timestamp 1681708930
transform 1 0 1532 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2517
timestamp 1681708930
transform 1 0 1476 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_2521
timestamp 1681708930
transform 1 0 1484 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_2518
timestamp 1681708930
transform 1 0 1508 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2486
timestamp 1681708930
transform 1 0 1588 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2522
timestamp 1681708930
transform 1 0 1532 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2598
timestamp 1681708930
transform 1 0 1444 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2599
timestamp 1681708930
transform 1 0 1452 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2559
timestamp 1681708930
transform 1 0 1452 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2577
timestamp 1681708930
transform 1 0 1412 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_2600
timestamp 1681708930
transform 1 0 1500 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2601
timestamp 1681708930
transform 1 0 1508 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2560
timestamp 1681708930
transform 1 0 1508 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2578
timestamp 1681708930
transform 1 0 1484 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2519
timestamp 1681708930
transform 1 0 1556 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2455
timestamp 1681708930
transform 1 0 1644 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_2523
timestamp 1681708930
transform 1 0 1588 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2602
timestamp 1681708930
transform 1 0 1556 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2603
timestamp 1681708930
transform 1 0 1564 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2579
timestamp 1681708930
transform 1 0 1540 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2520
timestamp 1681708930
transform 1 0 1612 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2487
timestamp 1681708930
transform 1 0 1668 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2488
timestamp 1681708930
transform 1 0 1700 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2524
timestamp 1681708930
transform 1 0 1636 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2525
timestamp 1681708930
transform 1 0 1644 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2604
timestamp 1681708930
transform 1 0 1612 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2526
timestamp 1681708930
transform 1 0 1700 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2605
timestamp 1681708930
transform 1 0 1668 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2606
timestamp 1681708930
transform 1 0 1676 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2580
timestamp 1681708930
transform 1 0 1620 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2581
timestamp 1681708930
transform 1 0 1644 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2418
timestamp 1681708930
transform 1 0 1748 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2419
timestamp 1681708930
transform 1 0 1772 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2420
timestamp 1681708930
transform 1 0 1820 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2489
timestamp 1681708930
transform 1 0 1788 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2527
timestamp 1681708930
transform 1 0 1788 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_2521
timestamp 1681708930
transform 1 0 1812 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2456
timestamp 1681708930
transform 1 0 1836 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2490
timestamp 1681708930
transform 1 0 1828 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2528
timestamp 1681708930
transform 1 0 1820 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2529
timestamp 1681708930
transform 1 0 1828 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2607
timestamp 1681708930
transform 1 0 1724 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2608
timestamp 1681708930
transform 1 0 1740 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2561
timestamp 1681708930
transform 1 0 1724 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2522
timestamp 1681708930
transform 1 0 1844 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_2530
timestamp 1681708930
transform 1 0 1852 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_2562
timestamp 1681708930
transform 1 0 1836 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2582
timestamp 1681708930
transform 1 0 1844 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2421
timestamp 1681708930
transform 1 0 1884 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2457
timestamp 1681708930
transform 1 0 1900 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2523
timestamp 1681708930
transform 1 0 1884 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_2531
timestamp 1681708930
transform 1 0 1892 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2609
timestamp 1681708930
transform 1 0 1876 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2610
timestamp 1681708930
transform 1 0 1884 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2611
timestamp 1681708930
transform 1 0 1900 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2524
timestamp 1681708930
transform 1 0 1916 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_2612
timestamp 1681708930
transform 1 0 1932 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2458
timestamp 1681708930
transform 1 0 1988 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2491
timestamp 1681708930
transform 1 0 1948 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2492
timestamp 1681708930
transform 1 0 1972 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2532
timestamp 1681708930
transform 1 0 1948 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2533
timestamp 1681708930
transform 1 0 1972 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_2459
timestamp 1681708930
transform 1 0 2004 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2434
timestamp 1681708930
transform 1 0 2020 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_2613
timestamp 1681708930
transform 1 0 2020 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2460
timestamp 1681708930
transform 1 0 2036 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2412
timestamp 1681708930
transform 1 0 2076 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2461
timestamp 1681708930
transform 1 0 2084 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2422
timestamp 1681708930
transform 1 0 2140 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2435
timestamp 1681708930
transform 1 0 2132 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2462
timestamp 1681708930
transform 1 0 2108 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2493
timestamp 1681708930
transform 1 0 2060 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2494
timestamp 1681708930
transform 1 0 2092 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2534
timestamp 1681708930
transform 1 0 2060 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2535
timestamp 1681708930
transform 1 0 2092 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2614
timestamp 1681708930
transform 1 0 2044 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2525
timestamp 1681708930
transform 1 0 2100 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_2536
timestamp 1681708930
transform 1 0 2116 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2537
timestamp 1681708930
transform 1 0 2132 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_2540
timestamp 1681708930
transform 1 0 2092 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2423
timestamp 1681708930
transform 1 0 2172 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2436
timestamp 1681708930
transform 1 0 2244 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2463
timestamp 1681708930
transform 1 0 2228 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2495
timestamp 1681708930
transform 1 0 2148 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2496
timestamp 1681708930
transform 1 0 2188 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2497
timestamp 1681708930
transform 1 0 2204 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2413
timestamp 1681708930
transform 1 0 2300 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2498
timestamp 1681708930
transform 1 0 2268 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2538
timestamp 1681708930
transform 1 0 2148 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2539
timestamp 1681708930
transform 1 0 2188 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2540
timestamp 1681708930
transform 1 0 2244 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2541
timestamp 1681708930
transform 1 0 2268 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2542
timestamp 1681708930
transform 1 0 2300 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2615
timestamp 1681708930
transform 1 0 2100 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2616
timestamp 1681708930
transform 1 0 2108 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2617
timestamp 1681708930
transform 1 0 2124 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2618
timestamp 1681708930
transform 1 0 2132 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2541
timestamp 1681708930
transform 1 0 2140 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_2619
timestamp 1681708930
transform 1 0 2164 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2620
timestamp 1681708930
transform 1 0 2300 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2414
timestamp 1681708930
transform 1 0 2372 0 1 1065
box -3 -3 3 3
use M2_M1  M2_M1_2469
timestamp 1681708930
transform 1 0 2356 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_2478
timestamp 1681708930
transform 1 0 2356 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2543
timestamp 1681708930
transform 1 0 2348 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2544
timestamp 1681708930
transform 1 0 2364 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_2415
timestamp 1681708930
transform 1 0 2396 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2526
timestamp 1681708930
transform 1 0 2388 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2542
timestamp 1681708930
transform 1 0 2364 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2543
timestamp 1681708930
transform 1 0 2380 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_2621
timestamp 1681708930
transform 1 0 2388 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2563
timestamp 1681708930
transform 1 0 2356 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_2636
timestamp 1681708930
transform 1 0 2380 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2479
timestamp 1681708930
transform 1 0 2428 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2480
timestamp 1681708930
transform 1 0 2460 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2481
timestamp 1681708930
transform 1 0 2476 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2545
timestamp 1681708930
transform 1 0 2444 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_2499
timestamp 1681708930
transform 1 0 2484 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2622
timestamp 1681708930
transform 1 0 2452 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2623
timestamp 1681708930
transform 1 0 2476 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2583
timestamp 1681708930
transform 1 0 2452 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_2470
timestamp 1681708930
transform 1 0 2508 0 1 1035
box -2 -2 2 2
use M3_M2  M3_M2_2527
timestamp 1681708930
transform 1 0 2508 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_2546
timestamp 1681708930
transform 1 0 2516 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2624
timestamp 1681708930
transform 1 0 2500 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2584
timestamp 1681708930
transform 1 0 2508 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2528
timestamp 1681708930
transform 1 0 2524 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_2625
timestamp 1681708930
transform 1 0 2540 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2564
timestamp 1681708930
transform 1 0 2540 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_2637
timestamp 1681708930
transform 1 0 2556 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_2464
timestamp 1681708930
transform 1 0 2564 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2465
timestamp 1681708930
transform 1 0 2580 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2466
timestamp 1681708930
transform 1 0 2596 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_2482
timestamp 1681708930
transform 1 0 2564 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_2500
timestamp 1681708930
transform 1 0 2580 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_2547
timestamp 1681708930
transform 1 0 2580 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2548
timestamp 1681708930
transform 1 0 2596 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_2585
timestamp 1681708930
transform 1 0 2564 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_2626
timestamp 1681708930
transform 1 0 2588 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2627
timestamp 1681708930
transform 1 0 2604 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2549
timestamp 1681708930
transform 1 0 2620 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2628
timestamp 1681708930
transform 1 0 2628 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_2586
timestamp 1681708930
transform 1 0 2620 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2529
timestamp 1681708930
transform 1 0 2644 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_2629
timestamp 1681708930
transform 1 0 2644 0 1 1005
box -2 -2 2 2
use top_mod_new_VIA0  top_mod_new_VIA0_32
timestamp 1681708930
transform 1 0 48 0 1 970
box -10 -3 10 3
use XNOR2X1  XNOR2X1_40
timestamp 1681708930
transform 1 0 72 0 1 970
box -8 -3 64 105
use NAND2X1  NAND2X1_59
timestamp 1681708930
transform 1 0 128 0 1 970
box -8 -3 32 105
use M3_M2  M3_M2_2587
timestamp 1681708930
transform 1 0 196 0 1 975
box -3 -3 3 3
use AOI22X1  AOI22X1_55
timestamp 1681708930
transform 1 0 152 0 1 970
box -8 -3 46 105
use INVX2  INVX2_166
timestamp 1681708930
transform 1 0 192 0 1 970
box -9 -3 26 105
use NOR2X1  NOR2X1_57
timestamp 1681708930
transform 1 0 208 0 1 970
box -8 -3 32 105
use M3_M2  M3_M2_2588
timestamp 1681708930
transform 1 0 252 0 1 975
box -3 -3 3 3
use OAI22X1  OAI22X1_23
timestamp 1681708930
transform 1 0 232 0 1 970
box -8 -3 46 105
use NAND3X1  NAND3X1_93
timestamp 1681708930
transform -1 0 304 0 1 970
box -8 -3 40 105
use NAND2X1  NAND2X1_60
timestamp 1681708930
transform 1 0 304 0 1 970
box -8 -3 32 105
use M3_M2  M3_M2_2589
timestamp 1681708930
transform 1 0 340 0 1 975
box -3 -3 3 3
use INVX2  INVX2_167
timestamp 1681708930
transform -1 0 344 0 1 970
box -9 -3 26 105
use FILL  FILL_1011
timestamp 1681708930
transform 1 0 344 0 1 970
box -8 -3 16 105
use FILL  FILL_1012
timestamp 1681708930
transform 1 0 352 0 1 970
box -8 -3 16 105
use INVX2  INVX2_168
timestamp 1681708930
transform -1 0 376 0 1 970
box -9 -3 26 105
use M3_M2  M3_M2_2590
timestamp 1681708930
transform 1 0 420 0 1 975
box -3 -3 3 3
use XOR2X1  XOR2X1_122
timestamp 1681708930
transform 1 0 376 0 1 970
box -8 -3 64 105
use OAI22X1  OAI22X1_24
timestamp 1681708930
transform 1 0 432 0 1 970
box -8 -3 46 105
use M3_M2  M3_M2_2591
timestamp 1681708930
transform 1 0 532 0 1 975
box -3 -3 3 3
use XOR2X1  XOR2X1_123
timestamp 1681708930
transform -1 0 528 0 1 970
box -8 -3 64 105
use FILL  FILL_1013
timestamp 1681708930
transform 1 0 528 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_2592
timestamp 1681708930
transform 1 0 572 0 1 975
box -3 -3 3 3
use AOI21X1  AOI21X1_36
timestamp 1681708930
transform -1 0 568 0 1 970
box -7 -3 39 105
use FILL  FILL_1014
timestamp 1681708930
transform 1 0 568 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_62
timestamp 1681708930
transform -1 0 608 0 1 970
box -8 -3 34 105
use INVX2  INVX2_169
timestamp 1681708930
transform -1 0 624 0 1 970
box -9 -3 26 105
use FILL  FILL_1015
timestamp 1681708930
transform 1 0 624 0 1 970
box -8 -3 16 105
use NOR2X1  NOR2X1_59
timestamp 1681708930
transform 1 0 632 0 1 970
box -8 -3 32 105
use AOI22X1  AOI22X1_56
timestamp 1681708930
transform 1 0 656 0 1 970
box -8 -3 46 105
use FILL  FILL_1023
timestamp 1681708930
transform 1 0 696 0 1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_61
timestamp 1681708930
transform -1 0 728 0 1 970
box -8 -3 32 105
use M3_M2  M3_M2_2593
timestamp 1681708930
transform 1 0 748 0 1 975
box -3 -3 3 3
use XOR2X1  XOR2X1_125
timestamp 1681708930
transform -1 0 784 0 1 970
box -8 -3 64 105
use XNOR2X1  XNOR2X1_41
timestamp 1681708930
transform -1 0 840 0 1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_126
timestamp 1681708930
transform 1 0 840 0 1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_127
timestamp 1681708930
transform -1 0 952 0 1 970
box -8 -3 64 105
use BUFX2  BUFX2_7
timestamp 1681708930
transform 1 0 952 0 1 970
box -5 -3 28 105
use XOR2X1  XOR2X1_128
timestamp 1681708930
transform 1 0 976 0 1 970
box -8 -3 64 105
use FILL  FILL_1024
timestamp 1681708930
transform 1 0 1032 0 1 970
box -8 -3 16 105
use FILL  FILL_1025
timestamp 1681708930
transform 1 0 1040 0 1 970
box -8 -3 16 105
use FILL  FILL_1042
timestamp 1681708930
transform 1 0 1048 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_64
timestamp 1681708930
transform -1 0 1088 0 1 970
box -8 -3 34 105
use FILL  FILL_1043
timestamp 1681708930
transform 1 0 1088 0 1 970
box -8 -3 16 105
use FILL  FILL_1044
timestamp 1681708930
transform 1 0 1096 0 1 970
box -8 -3 16 105
use FILL  FILL_1045
timestamp 1681708930
transform 1 0 1104 0 1 970
box -8 -3 16 105
use FILL  FILL_1046
timestamp 1681708930
transform 1 0 1112 0 1 970
box -8 -3 16 105
use FILL  FILL_1047
timestamp 1681708930
transform 1 0 1120 0 1 970
box -8 -3 16 105
use NOR2X1  NOR2X1_60
timestamp 1681708930
transform 1 0 1128 0 1 970
box -8 -3 32 105
use FILL  FILL_1048
timestamp 1681708930
transform 1 0 1152 0 1 970
box -8 -3 16 105
use FILL  FILL_1049
timestamp 1681708930
transform 1 0 1160 0 1 970
box -8 -3 16 105
use FILL  FILL_1050
timestamp 1681708930
transform 1 0 1168 0 1 970
box -8 -3 16 105
use FILL  FILL_1051
timestamp 1681708930
transform 1 0 1176 0 1 970
box -8 -3 16 105
use FILL  FILL_1058
timestamp 1681708930
transform 1 0 1184 0 1 970
box -8 -3 16 105
use INVX2  INVX2_172
timestamp 1681708930
transform 1 0 1192 0 1 970
box -9 -3 26 105
use FILL  FILL_1060
timestamp 1681708930
transform 1 0 1208 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_2594
timestamp 1681708930
transform 1 0 1228 0 1 975
box -3 -3 3 3
use FILL  FILL_1061
timestamp 1681708930
transform 1 0 1216 0 1 970
box -8 -3 16 105
use FILL  FILL_1062
timestamp 1681708930
transform 1 0 1224 0 1 970
box -8 -3 16 105
use FILL  FILL_1063
timestamp 1681708930
transform 1 0 1232 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_58
timestamp 1681708930
transform -1 0 1280 0 1 970
box -8 -3 46 105
use AOI21X1  AOI21X1_38
timestamp 1681708930
transform -1 0 1312 0 1 970
box -7 -3 39 105
use M3_M2  M3_M2_2595
timestamp 1681708930
transform 1 0 1324 0 1 975
box -3 -3 3 3
use NOR2X1  NOR2X1_61
timestamp 1681708930
transform 1 0 1312 0 1 970
box -8 -3 32 105
use XNOR2X1  XNOR2X1_42
timestamp 1681708930
transform -1 0 1392 0 1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_131
timestamp 1681708930
transform 1 0 1392 0 1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_132
timestamp 1681708930
transform 1 0 1448 0 1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_133
timestamp 1681708930
transform 1 0 1504 0 1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_134
timestamp 1681708930
transform 1 0 1560 0 1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_135
timestamp 1681708930
transform -1 0 1672 0 1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_136
timestamp 1681708930
transform 1 0 1672 0 1 970
box -8 -3 64 105
use DFFNEGX1  DFFNEGX1_67
timestamp 1681708930
transform 1 0 1728 0 1 970
box -8 -3 104 105
use FILL  FILL_1064
timestamp 1681708930
transform 1 0 1824 0 1 970
box -8 -3 16 105
use FILL  FILL_1078
timestamp 1681708930
transform 1 0 1832 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_2596
timestamp 1681708930
transform 1 0 1852 0 1 975
box -3 -3 3 3
use INVX2  INVX2_174
timestamp 1681708930
transform -1 0 1856 0 1 970
box -9 -3 26 105
use FILL  FILL_1079
timestamp 1681708930
transform 1 0 1856 0 1 970
box -8 -3 16 105
use FILL  FILL_1080
timestamp 1681708930
transform 1 0 1864 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_2597
timestamp 1681708930
transform 1 0 1892 0 1 975
box -3 -3 3 3
use AOI22X1  AOI22X1_60
timestamp 1681708930
transform -1 0 1912 0 1 970
box -8 -3 46 105
use FILL  FILL_1081
timestamp 1681708930
transform 1 0 1912 0 1 970
box -8 -3 16 105
use FILL  FILL_1086
timestamp 1681708930
transform 1 0 1920 0 1 970
box -8 -3 16 105
use FILL  FILL_1088
timestamp 1681708930
transform 1 0 1928 0 1 970
box -8 -3 16 105
use FILL  FILL_1090
timestamp 1681708930
transform 1 0 1936 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_2598
timestamp 1681708930
transform 1 0 2004 0 1 975
box -3 -3 3 3
use XOR2X1  XOR2X1_145
timestamp 1681708930
transform 1 0 1944 0 1 970
box -8 -3 64 105
use FILL  FILL_1091
timestamp 1681708930
transform 1 0 2000 0 1 970
box -8 -3 16 105
use FILL  FILL_1094
timestamp 1681708930
transform 1 0 2008 0 1 970
box -8 -3 16 105
use FILL  FILL_1095
timestamp 1681708930
transform 1 0 2016 0 1 970
box -8 -3 16 105
use FILL  FILL_1096
timestamp 1681708930
transform 1 0 2024 0 1 970
box -8 -3 16 105
use FILL  FILL_1097
timestamp 1681708930
transform 1 0 2032 0 1 970
box -8 -3 16 105
use XNOR2X1  XNOR2X1_43
timestamp 1681708930
transform -1 0 2096 0 1 970
box -8 -3 64 105
use AOI22X1  AOI22X1_61
timestamp 1681708930
transform 1 0 2096 0 1 970
box -8 -3 46 105
use INVX2  INVX2_175
timestamp 1681708930
transform 1 0 2136 0 1 970
box -9 -3 26 105
use M3_M2  M3_M2_2599
timestamp 1681708930
transform 1 0 2244 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_68
timestamp 1681708930
transform 1 0 2152 0 1 970
box -8 -3 104 105
use XOR2X1  XOR2X1_147
timestamp 1681708930
transform -1 0 2304 0 1 970
box -8 -3 64 105
use INVX2  INVX2_176
timestamp 1681708930
transform -1 0 2320 0 1 970
box -9 -3 26 105
use FILL  FILL_1098
timestamp 1681708930
transform 1 0 2320 0 1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_103
timestamp 1681708930
transform -1 0 2360 0 1 970
box -8 -3 40 105
use INVX2  INVX2_177
timestamp 1681708930
transform -1 0 2376 0 1 970
box -9 -3 26 105
use NOR2X1  NOR2X1_62
timestamp 1681708930
transform 1 0 2376 0 1 970
box -8 -3 32 105
use FILL  FILL_1099
timestamp 1681708930
transform 1 0 2400 0 1 970
box -8 -3 16 105
use FILL  FILL_1100
timestamp 1681708930
transform 1 0 2408 0 1 970
box -8 -3 16 105
use FILL  FILL_1117
timestamp 1681708930
transform 1 0 2416 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_2600
timestamp 1681708930
transform 1 0 2444 0 1 975
box -3 -3 3 3
use OAI21X1  OAI21X1_65
timestamp 1681708930
transform -1 0 2456 0 1 970
box -8 -3 34 105
use NAND3X1  NAND3X1_104
timestamp 1681708930
transform -1 0 2488 0 1 970
box -8 -3 40 105
use FILL  FILL_1118
timestamp 1681708930
transform 1 0 2488 0 1 970
box -8 -3 16 105
use FILL  FILL_1122
timestamp 1681708930
transform 1 0 2496 0 1 970
box -8 -3 16 105
use FILL  FILL_1124
timestamp 1681708930
transform 1 0 2504 0 1 970
box -8 -3 16 105
use NOR2X1  NOR2X1_64
timestamp 1681708930
transform -1 0 2536 0 1 970
box -8 -3 32 105
use FILL  FILL_1125
timestamp 1681708930
transform 1 0 2536 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_2601
timestamp 1681708930
transform 1 0 2556 0 1 975
box -3 -3 3 3
use FILL  FILL_1126
timestamp 1681708930
transform 1 0 2544 0 1 970
box -8 -3 16 105
use FILL  FILL_1127
timestamp 1681708930
transform 1 0 2552 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_66
timestamp 1681708930
transform -1 0 2592 0 1 970
box -8 -3 34 105
use INVX2  INVX2_179
timestamp 1681708930
transform -1 0 2608 0 1 970
box -9 -3 26 105
use FILL  FILL_1128
timestamp 1681708930
transform 1 0 2608 0 1 970
box -8 -3 16 105
use FILL  FILL_1129
timestamp 1681708930
transform 1 0 2616 0 1 970
box -8 -3 16 105
use FILL  FILL_1130
timestamp 1681708930
transform 1 0 2624 0 1 970
box -8 -3 16 105
use INVX2  INVX2_180
timestamp 1681708930
transform -1 0 2648 0 1 970
box -9 -3 26 105
use FILL  FILL_1131
timestamp 1681708930
transform 1 0 2648 0 1 970
box -8 -3 16 105
use FILL  FILL_1132
timestamp 1681708930
transform 1 0 2656 0 1 970
box -8 -3 16 105
use top_mod_new_VIA0  top_mod_new_VIA0_33
timestamp 1681708930
transform 1 0 2688 0 1 970
box -10 -3 10 3
use M2_M1  M2_M1_2646
timestamp 1681708930
transform 1 0 84 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_2668
timestamp 1681708930
transform 1 0 148 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2676
timestamp 1681708930
transform 1 0 84 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_2717
timestamp 1681708930
transform 1 0 108 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2718
timestamp 1681708930
transform 1 0 124 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2677
timestamp 1681708930
transform 1 0 156 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2618
timestamp 1681708930
transform 1 0 268 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2619
timestamp 1681708930
transform 1 0 300 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2620
timestamp 1681708930
transform 1 0 324 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2621
timestamp 1681708930
transform 1 0 340 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_2647
timestamp 1681708930
transform 1 0 252 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2648
timestamp 1681708930
transform 1 0 268 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2719
timestamp 1681708930
transform 1 0 164 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2720
timestamp 1681708930
transform 1 0 172 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2721
timestamp 1681708930
transform 1 0 228 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2695
timestamp 1681708930
transform 1 0 124 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2696
timestamp 1681708930
transform 1 0 172 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2697
timestamp 1681708930
transform 1 0 228 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2669
timestamp 1681708930
transform 1 0 276 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_2649
timestamp 1681708930
transform 1 0 316 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2722
timestamp 1681708930
transform 1 0 276 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2723
timestamp 1681708930
transform 1 0 292 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2698
timestamp 1681708930
transform 1 0 292 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2646
timestamp 1681708930
transform 1 0 372 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2650
timestamp 1681708930
transform 1 0 340 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2651
timestamp 1681708930
transform 1 0 364 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2773
timestamp 1681708930
transform 1 0 300 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2774
timestamp 1681708930
transform 1 0 324 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2775
timestamp 1681708930
transform 1 0 332 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_2622
timestamp 1681708930
transform 1 0 404 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2647
timestamp 1681708930
transform 1 0 412 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2652
timestamp 1681708930
transform 1 0 404 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2724
timestamp 1681708930
transform 1 0 372 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2725
timestamp 1681708930
transform 1 0 388 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2776
timestamp 1681708930
transform 1 0 364 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2793
timestamp 1681708930
transform 1 0 340 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_2794
timestamp 1681708930
transform 1 0 348 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_2734
timestamp 1681708930
transform 1 0 364 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2751
timestamp 1681708930
transform 1 0 348 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_2777
timestamp 1681708930
transform 1 0 396 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2795
timestamp 1681708930
transform 1 0 396 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_2735
timestamp 1681708930
transform 1 0 396 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2752
timestamp 1681708930
transform 1 0 380 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2602
timestamp 1681708930
transform 1 0 428 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_2653
timestamp 1681708930
transform 1 0 444 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2803
timestamp 1681708930
transform 1 0 428 0 1 895
box -2 -2 2 2
use M3_M2  M3_M2_2736
timestamp 1681708930
transform 1 0 436 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_2726
timestamp 1681708930
transform 1 0 460 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2623
timestamp 1681708930
transform 1 0 524 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2648
timestamp 1681708930
transform 1 0 516 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2649
timestamp 1681708930
transform 1 0 540 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2654
timestamp 1681708930
transform 1 0 516 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2655
timestamp 1681708930
transform 1 0 524 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2656
timestamp 1681708930
transform 1 0 540 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2727
timestamp 1681708930
transform 1 0 508 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2670
timestamp 1681708930
transform 1 0 548 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_2657
timestamp 1681708930
transform 1 0 564 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2658
timestamp 1681708930
transform 1 0 572 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2728
timestamp 1681708930
transform 1 0 548 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2678
timestamp 1681708930
transform 1 0 556 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_2729
timestamp 1681708930
transform 1 0 564 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2679
timestamp 1681708930
transform 1 0 572 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2603
timestamp 1681708930
transform 1 0 612 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2624
timestamp 1681708930
transform 1 0 596 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_2639
timestamp 1681708930
transform 1 0 588 0 1 945
box -2 -2 2 2
use M3_M2  M3_M2_2699
timestamp 1681708930
transform 1 0 580 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_2778
timestamp 1681708930
transform 1 0 588 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2796
timestamp 1681708930
transform 1 0 588 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_2730
timestamp 1681708930
transform 1 0 604 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2625
timestamp 1681708930
transform 1 0 628 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_2731
timestamp 1681708930
transform 1 0 628 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2779
timestamp 1681708930
transform 1 0 620 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_2718
timestamp 1681708930
transform 1 0 604 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2700
timestamp 1681708930
transform 1 0 628 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_2640
timestamp 1681708930
transform 1 0 660 0 1 945
box -2 -2 2 2
use M3_M2  M3_M2_2650
timestamp 1681708930
transform 1 0 684 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2659
timestamp 1681708930
transform 1 0 684 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_2701
timestamp 1681708930
transform 1 0 684 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2737
timestamp 1681708930
transform 1 0 676 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2626
timestamp 1681708930
transform 1 0 700 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_2660
timestamp 1681708930
transform 1 0 700 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2732
timestamp 1681708930
transform 1 0 700 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2627
timestamp 1681708930
transform 1 0 716 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_2733
timestamp 1681708930
transform 1 0 708 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2719
timestamp 1681708930
transform 1 0 700 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2651
timestamp 1681708930
transform 1 0 724 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2661
timestamp 1681708930
transform 1 0 724 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2734
timestamp 1681708930
transform 1 0 724 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2702
timestamp 1681708930
transform 1 0 724 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2628
timestamp 1681708930
transform 1 0 772 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_2641
timestamp 1681708930
transform 1 0 772 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2662
timestamp 1681708930
transform 1 0 764 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_2652
timestamp 1681708930
transform 1 0 788 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2780
timestamp 1681708930
transform 1 0 780 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_2738
timestamp 1681708930
transform 1 0 780 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2629
timestamp 1681708930
transform 1 0 812 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2653
timestamp 1681708930
transform 1 0 804 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2663
timestamp 1681708930
transform 1 0 812 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2781
timestamp 1681708930
transform 1 0 812 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2797
timestamp 1681708930
transform 1 0 804 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_2604
timestamp 1681708930
transform 1 0 828 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_2664
timestamp 1681708930
transform 1 0 844 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2735
timestamp 1681708930
transform 1 0 844 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2665
timestamp 1681708930
transform 1 0 892 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2666
timestamp 1681708930
transform 1 0 900 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_2605
timestamp 1681708930
transform 1 0 956 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2654
timestamp 1681708930
transform 1 0 948 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2667
timestamp 1681708930
transform 1 0 956 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2736
timestamp 1681708930
transform 1 0 916 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2737
timestamp 1681708930
transform 1 0 948 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2738
timestamp 1681708930
transform 1 0 964 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2655
timestamp 1681708930
transform 1 0 1012 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2739
timestamp 1681708930
transform 1 0 996 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2680
timestamp 1681708930
transform 1 0 1004 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2681
timestamp 1681708930
transform 1 0 1020 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_2740
timestamp 1681708930
transform 1 0 1028 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2782
timestamp 1681708930
transform 1 0 980 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_2703
timestamp 1681708930
transform 1 0 996 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_2783
timestamp 1681708930
transform 1 0 1004 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2784
timestamp 1681708930
transform 1 0 1012 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2798
timestamp 1681708930
transform 1 0 996 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_2720
timestamp 1681708930
transform 1 0 1004 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2671
timestamp 1681708930
transform 1 0 1052 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_2668
timestamp 1681708930
transform 1 0 1068 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2799
timestamp 1681708930
transform 1 0 1060 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_2739
timestamp 1681708930
transform 1 0 1060 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2672
timestamp 1681708930
transform 1 0 1076 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2656
timestamp 1681708930
transform 1 0 1100 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2669
timestamp 1681708930
transform 1 0 1100 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2670
timestamp 1681708930
transform 1 0 1116 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2671
timestamp 1681708930
transform 1 0 1124 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2741
timestamp 1681708930
transform 1 0 1108 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2704
timestamp 1681708930
transform 1 0 1108 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_2785
timestamp 1681708930
transform 1 0 1132 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2672
timestamp 1681708930
transform 1 0 1156 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2800
timestamp 1681708930
transform 1 0 1148 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_2673
timestamp 1681708930
transform 1 0 1180 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2786
timestamp 1681708930
transform 1 0 1172 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_2721
timestamp 1681708930
transform 1 0 1172 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_2674
timestamp 1681708930
transform 1 0 1196 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_2682
timestamp 1681708930
transform 1 0 1196 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2606
timestamp 1681708930
transform 1 0 1244 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2657
timestamp 1681708930
transform 1 0 1228 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2675
timestamp 1681708930
transform 1 0 1228 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2676
timestamp 1681708930
transform 1 0 1236 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2677
timestamp 1681708930
transform 1 0 1260 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2742
timestamp 1681708930
transform 1 0 1204 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2743
timestamp 1681708930
transform 1 0 1220 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2744
timestamp 1681708930
transform 1 0 1236 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2745
timestamp 1681708930
transform 1 0 1244 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2722
timestamp 1681708930
transform 1 0 1188 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2705
timestamp 1681708930
transform 1 0 1244 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2723
timestamp 1681708930
transform 1 0 1228 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2724
timestamp 1681708930
transform 1 0 1244 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2740
timestamp 1681708930
transform 1 0 1220 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2741
timestamp 1681708930
transform 1 0 1236 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2607
timestamp 1681708930
transform 1 0 1284 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2630
timestamp 1681708930
transform 1 0 1276 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_2642
timestamp 1681708930
transform 1 0 1276 0 1 945
box -2 -2 2 2
use M3_M2  M3_M2_2742
timestamp 1681708930
transform 1 0 1268 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2658
timestamp 1681708930
transform 1 0 1292 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2678
timestamp 1681708930
transform 1 0 1292 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_2631
timestamp 1681708930
transform 1 0 1316 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2683
timestamp 1681708930
transform 1 0 1308 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_2787
timestamp 1681708930
transform 1 0 1308 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_2632
timestamp 1681708930
transform 1 0 1356 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2659
timestamp 1681708930
transform 1 0 1332 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2679
timestamp 1681708930
transform 1 0 1332 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_2673
timestamp 1681708930
transform 1 0 1340 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2660
timestamp 1681708930
transform 1 0 1372 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2680
timestamp 1681708930
transform 1 0 1356 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2681
timestamp 1681708930
transform 1 0 1372 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_2684
timestamp 1681708930
transform 1 0 1348 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_2788
timestamp 1681708930
transform 1 0 1340 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2789
timestamp 1681708930
transform 1 0 1356 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_2743
timestamp 1681708930
transform 1 0 1324 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_2801
timestamp 1681708930
transform 1 0 1348 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_2725
timestamp 1681708930
transform 1 0 1356 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2608
timestamp 1681708930
transform 1 0 1444 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_2682
timestamp 1681708930
transform 1 0 1428 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2746
timestamp 1681708930
transform 1 0 1388 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2685
timestamp 1681708930
transform 1 0 1396 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2686
timestamp 1681708930
transform 1 0 1428 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2633
timestamp 1681708930
transform 1 0 1476 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2634
timestamp 1681708930
transform 1 0 1500 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_2683
timestamp 1681708930
transform 1 0 1484 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2684
timestamp 1681708930
transform 1 0 1532 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2685
timestamp 1681708930
transform 1 0 1540 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2747
timestamp 1681708930
transform 1 0 1452 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2748
timestamp 1681708930
transform 1 0 1484 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2749
timestamp 1681708930
transform 1 0 1508 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2726
timestamp 1681708930
transform 1 0 1412 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2706
timestamp 1681708930
transform 1 0 1444 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2744
timestamp 1681708930
transform 1 0 1428 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2753
timestamp 1681708930
transform 1 0 1388 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2707
timestamp 1681708930
transform 1 0 1508 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2745
timestamp 1681708930
transform 1 0 1484 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2635
timestamp 1681708930
transform 1 0 1668 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2636
timestamp 1681708930
transform 1 0 1700 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2661
timestamp 1681708930
transform 1 0 1644 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2686
timestamp 1681708930
transform 1 0 1644 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2687
timestamp 1681708930
transform 1 0 1652 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_2662
timestamp 1681708930
transform 1 0 1708 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2688
timestamp 1681708930
transform 1 0 1700 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2689
timestamp 1681708930
transform 1 0 1708 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2750
timestamp 1681708930
transform 1 0 1564 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2751
timestamp 1681708930
transform 1 0 1588 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2752
timestamp 1681708930
transform 1 0 1596 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2753
timestamp 1681708930
transform 1 0 1620 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2754
timestamp 1681708930
transform 1 0 1644 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2746
timestamp 1681708930
transform 1 0 1564 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2754
timestamp 1681708930
transform 1 0 1548 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2755
timestamp 1681708930
transform 1 0 1588 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2687
timestamp 1681708930
transform 1 0 1668 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2708
timestamp 1681708930
transform 1 0 1652 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_2690
timestamp 1681708930
transform 1 0 1756 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2755
timestamp 1681708930
transform 1 0 1732 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2709
timestamp 1681708930
transform 1 0 1708 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2710
timestamp 1681708930
transform 1 0 1732 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2747
timestamp 1681708930
transform 1 0 1724 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2748
timestamp 1681708930
transform 1 0 1780 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2609
timestamp 1681708930
transform 1 0 1796 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_2691
timestamp 1681708930
transform 1 0 1820 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2692
timestamp 1681708930
transform 1 0 1844 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2756
timestamp 1681708930
transform 1 0 1868 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2610
timestamp 1681708930
transform 1 0 1900 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2663
timestamp 1681708930
transform 1 0 1916 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2693
timestamp 1681708930
transform 1 0 1908 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2694
timestamp 1681708930
transform 1 0 1932 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_2688
timestamp 1681708930
transform 1 0 1932 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2749
timestamp 1681708930
transform 1 0 1932 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_2757
timestamp 1681708930
transform 1 0 1964 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2695
timestamp 1681708930
transform 1 0 1996 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_2637
timestamp 1681708930
transform 1 0 2036 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_2696
timestamp 1681708930
transform 1 0 2012 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_2638
timestamp 1681708930
transform 1 0 2076 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2664
timestamp 1681708930
transform 1 0 2068 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2697
timestamp 1681708930
transform 1 0 2060 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2698
timestamp 1681708930
transform 1 0 2068 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_2689
timestamp 1681708930
transform 1 0 2044 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2690
timestamp 1681708930
transform 1 0 2076 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2611
timestamp 1681708930
transform 1 0 2108 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2639
timestamp 1681708930
transform 1 0 2116 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2756
timestamp 1681708930
transform 1 0 2108 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2612
timestamp 1681708930
transform 1 0 2156 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2640
timestamp 1681708930
transform 1 0 2132 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_2699
timestamp 1681708930
transform 1 0 2124 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2700
timestamp 1681708930
transform 1 0 2156 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2758
timestamp 1681708930
transform 1 0 2124 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2759
timestamp 1681708930
transform 1 0 2132 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2760
timestamp 1681708930
transform 1 0 2148 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2757
timestamp 1681708930
transform 1 0 2148 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2613
timestamp 1681708930
transform 1 0 2172 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_2701
timestamp 1681708930
transform 1 0 2172 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_2727
timestamp 1681708930
transform 1 0 2172 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2641
timestamp 1681708930
transform 1 0 2228 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_2643
timestamp 1681708930
transform 1 0 2244 0 1 945
box -2 -2 2 2
use M3_M2  M3_M2_2665
timestamp 1681708930
transform 1 0 2252 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2644
timestamp 1681708930
transform 1 0 2260 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2702
timestamp 1681708930
transform 1 0 2236 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_2674
timestamp 1681708930
transform 1 0 2244 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_2761
timestamp 1681708930
transform 1 0 2188 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2762
timestamp 1681708930
transform 1 0 2212 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2711
timestamp 1681708930
transform 1 0 2188 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2712
timestamp 1681708930
transform 1 0 2212 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2758
timestamp 1681708930
transform 1 0 2196 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_2703
timestamp 1681708930
transform 1 0 2268 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2763
timestamp 1681708930
transform 1 0 2260 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2759
timestamp 1681708930
transform 1 0 2252 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_2704
timestamp 1681708930
transform 1 0 2276 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2764
timestamp 1681708930
transform 1 0 2284 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2713
timestamp 1681708930
transform 1 0 2284 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2642
timestamp 1681708930
transform 1 0 2308 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2666
timestamp 1681708930
transform 1 0 2300 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2705
timestamp 1681708930
transform 1 0 2300 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_2643
timestamp 1681708930
transform 1 0 2340 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2667
timestamp 1681708930
transform 1 0 2364 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_2706
timestamp 1681708930
transform 1 0 2364 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2765
timestamp 1681708930
transform 1 0 2332 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2714
timestamp 1681708930
transform 1 0 2364 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2728
timestamp 1681708930
transform 1 0 2332 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2729
timestamp 1681708930
transform 1 0 2356 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2644
timestamp 1681708930
transform 1 0 2380 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_2645
timestamp 1681708930
transform 1 0 2380 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2707
timestamp 1681708930
transform 1 0 2380 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_2691
timestamp 1681708930
transform 1 0 2388 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2715
timestamp 1681708930
transform 1 0 2396 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_2708
timestamp 1681708930
transform 1 0 2412 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_2730
timestamp 1681708930
transform 1 0 2412 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2645
timestamp 1681708930
transform 1 0 2428 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2614
timestamp 1681708930
transform 1 0 2476 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_2709
timestamp 1681708930
transform 1 0 2436 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_2692
timestamp 1681708930
transform 1 0 2436 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_2710
timestamp 1681708930
transform 1 0 2484 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2766
timestamp 1681708930
transform 1 0 2484 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_2731
timestamp 1681708930
transform 1 0 2468 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2693
timestamp 1681708930
transform 1 0 2500 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2615
timestamp 1681708930
transform 1 0 2516 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2616
timestamp 1681708930
transform 1 0 2540 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2617
timestamp 1681708930
transform 1 0 2604 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_2711
timestamp 1681708930
transform 1 0 2540 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2712
timestamp 1681708930
transform 1 0 2548 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2713
timestamp 1681708930
transform 1 0 2564 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2714
timestamp 1681708930
transform 1 0 2572 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2715
timestamp 1681708930
transform 1 0 2580 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2767
timestamp 1681708930
transform 1 0 2516 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2768
timestamp 1681708930
transform 1 0 2540 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2769
timestamp 1681708930
transform 1 0 2556 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2790
timestamp 1681708930
transform 1 0 2508 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2802
timestamp 1681708930
transform 1 0 2500 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_2760
timestamp 1681708930
transform 1 0 2500 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2716
timestamp 1681708930
transform 1 0 2516 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_2791
timestamp 1681708930
transform 1 0 2532 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_2717
timestamp 1681708930
transform 1 0 2548 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2675
timestamp 1681708930
transform 1 0 2596 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_2716
timestamp 1681708930
transform 1 0 2604 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2770
timestamp 1681708930
transform 1 0 2596 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2771
timestamp 1681708930
transform 1 0 2604 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2792
timestamp 1681708930
transform 1 0 2580 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_2732
timestamp 1681708930
transform 1 0 2532 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2750
timestamp 1681708930
transform 1 0 2516 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2761
timestamp 1681708930
transform 1 0 2524 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2733
timestamp 1681708930
transform 1 0 2580 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2694
timestamp 1681708930
transform 1 0 2636 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_2772
timestamp 1681708930
transform 1 0 2644 0 1 925
box -2 -2 2 2
use top_mod_new_VIA0  top_mod_new_VIA0_34
timestamp 1681708930
transform 1 0 24 0 1 870
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_65
timestamp 1681708930
transform 1 0 72 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_66
timestamp 1681708930
transform -1 0 264 0 -1 970
box -8 -3 104 105
use OAI21X1  OAI21X1_63
timestamp 1681708930
transform 1 0 264 0 -1 970
box -8 -3 34 105
use NAND3X1  NAND3X1_94
timestamp 1681708930
transform -1 0 328 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_95
timestamp 1681708930
transform 1 0 328 0 -1 970
box -8 -3 40 105
use AND2X2  AND2X2_3
timestamp 1681708930
transform 1 0 360 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_96
timestamp 1681708930
transform 1 0 392 0 -1 970
box -8 -3 40 105
use FILL  FILL_1016
timestamp 1681708930
transform 1 0 424 0 -1 970
box -8 -3 16 105
use FILL  FILL_1017
timestamp 1681708930
transform 1 0 432 0 -1 970
box -8 -3 16 105
use XOR2X1  XOR2X1_124
timestamp 1681708930
transform -1 0 496 0 -1 970
box -8 -3 64 105
use FILL  FILL_1018
timestamp 1681708930
transform 1 0 496 0 -1 970
box -8 -3 16 105
use FILL  FILL_1019
timestamp 1681708930
transform 1 0 504 0 -1 970
box -8 -3 16 105
use FILL  FILL_1020
timestamp 1681708930
transform 1 0 512 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_25
timestamp 1681708930
transform 1 0 520 0 -1 970
box -8 -3 46 105
use NOR2X1  NOR2X1_58
timestamp 1681708930
transform -1 0 584 0 -1 970
box -8 -3 32 105
use FILL  FILL_1021
timestamp 1681708930
transform 1 0 584 0 -1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_97
timestamp 1681708930
transform 1 0 592 0 -1 970
box -8 -3 40 105
use FILL  FILL_1022
timestamp 1681708930
transform 1 0 624 0 -1 970
box -8 -3 16 105
use FILL  FILL_1026
timestamp 1681708930
transform 1 0 632 0 -1 970
box -8 -3 16 105
use FILL  FILL_1027
timestamp 1681708930
transform 1 0 640 0 -1 970
box -8 -3 16 105
use FILL  FILL_1028
timestamp 1681708930
transform 1 0 648 0 -1 970
box -8 -3 16 105
use FILL  FILL_1029
timestamp 1681708930
transform 1 0 656 0 -1 970
box -8 -3 16 105
use AOI21X1  AOI21X1_37
timestamp 1681708930
transform -1 0 696 0 -1 970
box -7 -3 39 105
use FILL  FILL_1030
timestamp 1681708930
transform 1 0 696 0 -1 970
box -8 -3 16 105
use FILL  FILL_1031
timestamp 1681708930
transform 1 0 704 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_170
timestamp 1681708930
transform -1 0 728 0 -1 970
box -9 -3 26 105
use FILL  FILL_1032
timestamp 1681708930
transform 1 0 728 0 -1 970
box -8 -3 16 105
use FILL  FILL_1033
timestamp 1681708930
transform 1 0 736 0 -1 970
box -8 -3 16 105
use OR2X1  OR2X1_17
timestamp 1681708930
transform -1 0 776 0 -1 970
box -8 -3 40 105
use FILL  FILL_1034
timestamp 1681708930
transform 1 0 776 0 -1 970
box -8 -3 16 105
use FILL  FILL_1035
timestamp 1681708930
transform 1 0 784 0 -1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_98
timestamp 1681708930
transform -1 0 824 0 -1 970
box -8 -3 40 105
use FILL  FILL_1036
timestamp 1681708930
transform 1 0 824 0 -1 970
box -8 -3 16 105
use FILL  FILL_1037
timestamp 1681708930
transform 1 0 832 0 -1 970
box -8 -3 16 105
use XOR2X1  XOR2X1_129
timestamp 1681708930
transform -1 0 896 0 -1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_130
timestamp 1681708930
transform -1 0 952 0 -1 970
box -8 -3 64 105
use FILL  FILL_1038
timestamp 1681708930
transform 1 0 952 0 -1 970
box -8 -3 16 105
use FILL  FILL_1039
timestamp 1681708930
transform 1 0 960 0 -1 970
box -8 -3 16 105
use FILL  FILL_1040
timestamp 1681708930
transform 1 0 968 0 -1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_99
timestamp 1681708930
transform -1 0 1008 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_100
timestamp 1681708930
transform -1 0 1040 0 -1 970
box -8 -3 40 105
use FILL  FILL_1041
timestamp 1681708930
transform 1 0 1040 0 -1 970
box -8 -3 16 105
use FILL  FILL_1052
timestamp 1681708930
transform 1 0 1048 0 -1 970
box -8 -3 16 105
use FILL  FILL_1053
timestamp 1681708930
transform 1 0 1056 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_171
timestamp 1681708930
transform 1 0 1064 0 -1 970
box -9 -3 26 105
use FILL  FILL_1054
timestamp 1681708930
transform 1 0 1080 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_57
timestamp 1681708930
transform -1 0 1128 0 -1 970
box -8 -3 46 105
use FILL  FILL_1055
timestamp 1681708930
transform 1 0 1128 0 -1 970
box -8 -3 16 105
use FILL  FILL_1056
timestamp 1681708930
transform 1 0 1136 0 -1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_101
timestamp 1681708930
transform 1 0 1144 0 -1 970
box -8 -3 40 105
use FILL  FILL_1057
timestamp 1681708930
transform 1 0 1176 0 -1 970
box -8 -3 16 105
use FILL  FILL_1059
timestamp 1681708930
transform 1 0 1184 0 -1 970
box -8 -3 16 105
use FILL  FILL_1065
timestamp 1681708930
transform 1 0 1192 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_59
timestamp 1681708930
transform -1 0 1240 0 -1 970
box -8 -3 46 105
use OR2X1  OR2X1_18
timestamp 1681708930
transform -1 0 1272 0 -1 970
box -8 -3 40 105
use FILL  FILL_1066
timestamp 1681708930
transform 1 0 1272 0 -1 970
box -8 -3 16 105
use FILL  FILL_1067
timestamp 1681708930
transform 1 0 1280 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_62
timestamp 1681708930
transform 1 0 1288 0 -1 970
box -8 -3 32 105
use FILL  FILL_1068
timestamp 1681708930
transform 1 0 1312 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_173
timestamp 1681708930
transform -1 0 1336 0 -1 970
box -9 -3 26 105
use NAND3X1  NAND3X1_102
timestamp 1681708930
transform -1 0 1368 0 -1 970
box -8 -3 40 105
use XOR2X1  XOR2X1_137
timestamp 1681708930
transform -1 0 1424 0 -1 970
box -8 -3 64 105
use M3_M2  M3_M2_2762
timestamp 1681708930
transform 1 0 1452 0 1 875
box -3 -3 3 3
use XOR2X1  XOR2X1_138
timestamp 1681708930
transform 1 0 1424 0 -1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_139
timestamp 1681708930
transform 1 0 1480 0 -1 970
box -8 -3 64 105
use M3_M2  M3_M2_2763
timestamp 1681708930
transform 1 0 1596 0 1 875
box -3 -3 3 3
use XOR2X1  XOR2X1_140
timestamp 1681708930
transform 1 0 1536 0 -1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_141
timestamp 1681708930
transform -1 0 1648 0 -1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_142
timestamp 1681708930
transform -1 0 1704 0 -1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_143
timestamp 1681708930
transform 1 0 1704 0 -1 970
box -8 -3 64 105
use FILL  FILL_1069
timestamp 1681708930
transform 1 0 1760 0 -1 970
box -8 -3 16 105
use FILL  FILL_1070
timestamp 1681708930
transform 1 0 1768 0 -1 970
box -8 -3 16 105
use FILL  FILL_1071
timestamp 1681708930
transform 1 0 1776 0 -1 970
box -8 -3 16 105
use FILL  FILL_1072
timestamp 1681708930
transform 1 0 1784 0 -1 970
box -8 -3 16 105
use FILL  FILL_1073
timestamp 1681708930
transform 1 0 1792 0 -1 970
box -8 -3 16 105
use FILL  FILL_1074
timestamp 1681708930
transform 1 0 1800 0 -1 970
box -8 -3 16 105
use FILL  FILL_1075
timestamp 1681708930
transform 1 0 1808 0 -1 970
box -8 -3 16 105
use FILL  FILL_1076
timestamp 1681708930
transform 1 0 1816 0 -1 970
box -8 -3 16 105
use FILL  FILL_1077
timestamp 1681708930
transform 1 0 1824 0 -1 970
box -8 -3 16 105
use FILL  FILL_1082
timestamp 1681708930
transform 1 0 1832 0 -1 970
box -8 -3 16 105
use XOR2X1  XOR2X1_144
timestamp 1681708930
transform 1 0 1840 0 -1 970
box -8 -3 64 105
use FILL  FILL_1083
timestamp 1681708930
transform 1 0 1896 0 -1 970
box -8 -3 16 105
use FILL  FILL_1084
timestamp 1681708930
transform 1 0 1904 0 -1 970
box -8 -3 16 105
use FILL  FILL_1085
timestamp 1681708930
transform 1 0 1912 0 -1 970
box -8 -3 16 105
use FILL  FILL_1087
timestamp 1681708930
transform 1 0 1920 0 -1 970
box -8 -3 16 105
use FILL  FILL_1089
timestamp 1681708930
transform 1 0 1928 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_2764
timestamp 1681708930
transform 1 0 1956 0 1 875
box -3 -3 3 3
use XOR2X1  XOR2X1_146
timestamp 1681708930
transform 1 0 1936 0 -1 970
box -8 -3 64 105
use FILL  FILL_1092
timestamp 1681708930
transform 1 0 1992 0 -1 970
box -8 -3 16 105
use FILL  FILL_1093
timestamp 1681708930
transform 1 0 2000 0 -1 970
box -8 -3 16 105
use XOR2X1  XOR2X1_148
timestamp 1681708930
transform 1 0 2008 0 -1 970
box -8 -3 64 105
use FILL  FILL_1101
timestamp 1681708930
transform 1 0 2064 0 -1 970
box -8 -3 16 105
use FILL  FILL_1102
timestamp 1681708930
transform 1 0 2072 0 -1 970
box -8 -3 16 105
use FILL  FILL_1103
timestamp 1681708930
transform 1 0 2080 0 -1 970
box -8 -3 16 105
use FILL  FILL_1104
timestamp 1681708930
transform 1 0 2088 0 -1 970
box -8 -3 16 105
use FILL  FILL_1105
timestamp 1681708930
transform 1 0 2096 0 -1 970
box -8 -3 16 105
use FILL  FILL_1106
timestamp 1681708930
transform 1 0 2104 0 -1 970
box -8 -3 16 105
use FILL  FILL_1107
timestamp 1681708930
transform 1 0 2112 0 -1 970
box -8 -3 16 105
use FILL  FILL_1108
timestamp 1681708930
transform 1 0 2120 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_62
timestamp 1681708930
transform -1 0 2168 0 -1 970
box -8 -3 46 105
use FILL  FILL_1109
timestamp 1681708930
transform 1 0 2168 0 -1 970
box -8 -3 16 105
use FILL  FILL_1110
timestamp 1681708930
transform 1 0 2176 0 -1 970
box -8 -3 16 105
use XOR2X1  XOR2X1_149
timestamp 1681708930
transform 1 0 2184 0 -1 970
box -8 -3 64 105
use NOR2X1  NOR2X1_63
timestamp 1681708930
transform 1 0 2240 0 -1 970
box -8 -3 32 105
use FILL  FILL_1111
timestamp 1681708930
transform 1 0 2264 0 -1 970
box -8 -3 16 105
use FILL  FILL_1112
timestamp 1681708930
transform 1 0 2272 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_178
timestamp 1681708930
transform 1 0 2280 0 -1 970
box -9 -3 26 105
use FILL  FILL_1113
timestamp 1681708930
transform 1 0 2296 0 -1 970
box -8 -3 16 105
use FILL  FILL_1114
timestamp 1681708930
transform 1 0 2304 0 -1 970
box -8 -3 16 105
use XNOR2X1  XNOR2X1_44
timestamp 1681708930
transform -1 0 2368 0 -1 970
box -8 -3 64 105
use FILL  FILL_1115
timestamp 1681708930
transform 1 0 2368 0 -1 970
box -8 -3 16 105
use AOI21X1  AOI21X1_39
timestamp 1681708930
transform -1 0 2408 0 -1 970
box -7 -3 39 105
use FILL  FILL_1116
timestamp 1681708930
transform 1 0 2408 0 -1 970
box -8 -3 16 105
use FILL  FILL_1119
timestamp 1681708930
transform 1 0 2416 0 -1 970
box -8 -3 16 105
use FILL  FILL_1120
timestamp 1681708930
transform 1 0 2424 0 -1 970
box -8 -3 16 105
use XNOR2X1  XNOR2X1_45
timestamp 1681708930
transform -1 0 2488 0 -1 970
box -8 -3 64 105
use FILL  FILL_1121
timestamp 1681708930
transform 1 0 2488 0 -1 970
box -8 -3 16 105
use FILL  FILL_1123
timestamp 1681708930
transform 1 0 2496 0 -1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_105
timestamp 1681708930
transform 1 0 2504 0 -1 970
box -8 -3 40 105
use AOI22X1  AOI22X1_63
timestamp 1681708930
transform -1 0 2576 0 -1 970
box -8 -3 46 105
use OAI21X1  OAI21X1_67
timestamp 1681708930
transform -1 0 2608 0 -1 970
box -8 -3 34 105
use XNOR2X1  XNOR2X1_46
timestamp 1681708930
transform 1 0 2608 0 -1 970
box -8 -3 64 105
use top_mod_new_VIA0  top_mod_new_VIA0_35
timestamp 1681708930
transform 1 0 2712 0 1 870
box -10 -3 10 3
use M3_M2  M3_M2_2788
timestamp 1681708930
transform 1 0 188 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_2810
timestamp 1681708930
transform 1 0 188 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2833
timestamp 1681708930
transform 1 0 76 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2840
timestamp 1681708930
transform 1 0 84 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_2834
timestamp 1681708930
transform 1 0 132 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2841
timestamp 1681708930
transform 1 0 172 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_2915
timestamp 1681708930
transform 1 0 156 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2916
timestamp 1681708930
transform 1 0 172 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2917
timestamp 1681708930
transform 1 0 188 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2874
timestamp 1681708930
transform 1 0 132 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2804
timestamp 1681708930
transform 1 0 220 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2835
timestamp 1681708930
transform 1 0 212 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2875
timestamp 1681708930
transform 1 0 188 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2789
timestamp 1681708930
transform 1 0 324 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_2836
timestamp 1681708930
transform 1 0 284 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2837
timestamp 1681708930
transform 1 0 316 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2838
timestamp 1681708930
transform 1 0 324 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2918
timestamp 1681708930
transform 1 0 220 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2919
timestamp 1681708930
transform 1 0 236 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2861
timestamp 1681708930
transform 1 0 284 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2805
timestamp 1681708930
transform 1 0 348 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2806
timestamp 1681708930
transform 1 0 364 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2839
timestamp 1681708930
transform 1 0 348 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2840
timestamp 1681708930
transform 1 0 364 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2862
timestamp 1681708930
transform 1 0 348 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_2920
timestamp 1681708930
transform 1 0 356 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2841
timestamp 1681708930
transform 1 0 380 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2921
timestamp 1681708930
transform 1 0 372 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2807
timestamp 1681708930
transform 1 0 388 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2842
timestamp 1681708930
transform 1 0 388 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2922
timestamp 1681708930
transform 1 0 396 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2808
timestamp 1681708930
transform 1 0 420 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2843
timestamp 1681708930
transform 1 0 404 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2844
timestamp 1681708930
transform 1 0 420 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2863
timestamp 1681708930
transform 1 0 404 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_2923
timestamp 1681708930
transform 1 0 428 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2924
timestamp 1681708930
transform 1 0 436 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2876
timestamp 1681708930
transform 1 0 428 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_2845
timestamp 1681708930
transform 1 0 444 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2877
timestamp 1681708930
transform 1 0 452 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2864
timestamp 1681708930
transform 1 0 484 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2790
timestamp 1681708930
transform 1 0 500 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_2846
timestamp 1681708930
transform 1 0 508 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2925
timestamp 1681708930
transform 1 0 500 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2811
timestamp 1681708930
transform 1 0 524 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_2780
timestamp 1681708930
transform 1 0 564 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2791
timestamp 1681708930
transform 1 0 564 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2809
timestamp 1681708930
transform 1 0 564 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2847
timestamp 1681708930
transform 1 0 564 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2810
timestamp 1681708930
transform 1 0 588 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2848
timestamp 1681708930
transform 1 0 580 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2849
timestamp 1681708930
transform 1 0 596 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2926
timestamp 1681708930
transform 1 0 572 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2927
timestamp 1681708930
transform 1 0 612 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2878
timestamp 1681708930
transform 1 0 612 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2897
timestamp 1681708930
transform 1 0 604 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_2850
timestamp 1681708930
transform 1 0 636 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2811
timestamp 1681708930
transform 1 0 644 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2928
timestamp 1681708930
transform 1 0 644 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2879
timestamp 1681708930
transform 1 0 644 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2781
timestamp 1681708930
transform 1 0 668 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2792
timestamp 1681708930
transform 1 0 668 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_2804
timestamp 1681708930
transform 1 0 692 0 1 835
box -2 -2 2 2
use M3_M2  M3_M2_2793
timestamp 1681708930
transform 1 0 708 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_2812
timestamp 1681708930
transform 1 0 676 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2851
timestamp 1681708930
transform 1 0 668 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2812
timestamp 1681708930
transform 1 0 692 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2782
timestamp 1681708930
transform 1 0 740 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_2813
timestamp 1681708930
transform 1 0 700 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_2813
timestamp 1681708930
transform 1 0 724 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2852
timestamp 1681708930
transform 1 0 684 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2853
timestamp 1681708930
transform 1 0 708 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2854
timestamp 1681708930
transform 1 0 724 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2855
timestamp 1681708930
transform 1 0 740 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2929
timestamp 1681708930
transform 1 0 684 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2880
timestamp 1681708930
transform 1 0 676 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2898
timestamp 1681708930
transform 1 0 684 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_2930
timestamp 1681708930
transform 1 0 716 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2865
timestamp 1681708930
transform 1 0 724 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_2931
timestamp 1681708930
transform 1 0 732 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2773
timestamp 1681708930
transform 1 0 764 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_2856
timestamp 1681708930
transform 1 0 756 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2783
timestamp 1681708930
transform 1 0 812 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2794
timestamp 1681708930
transform 1 0 788 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2795
timestamp 1681708930
transform 1 0 812 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2814
timestamp 1681708930
transform 1 0 796 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2814
timestamp 1681708930
transform 1 0 820 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2932
timestamp 1681708930
transform 1 0 764 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2842
timestamp 1681708930
transform 1 0 820 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_2857
timestamp 1681708930
transform 1 0 836 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2899
timestamp 1681708930
transform 1 0 772 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_2933
timestamp 1681708930
transform 1 0 860 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2934
timestamp 1681708930
transform 1 0 868 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2796
timestamp 1681708930
transform 1 0 892 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_2815
timestamp 1681708930
transform 1 0 908 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2858
timestamp 1681708930
transform 1 0 900 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2866
timestamp 1681708930
transform 1 0 900 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_2805
timestamp 1681708930
transform 1 0 932 0 1 835
box -2 -2 2 2
use M3_M2  M3_M2_2797
timestamp 1681708930
transform 1 0 940 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2815
timestamp 1681708930
transform 1 0 924 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2816
timestamp 1681708930
transform 1 0 940 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2859
timestamp 1681708930
transform 1 0 924 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2806
timestamp 1681708930
transform 1 0 964 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_2817
timestamp 1681708930
transform 1 0 956 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_2816
timestamp 1681708930
transform 1 0 972 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2818
timestamp 1681708930
transform 1 0 980 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2860
timestamp 1681708930
transform 1 0 972 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2861
timestamp 1681708930
transform 1 0 988 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2867
timestamp 1681708930
transform 1 0 988 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2774
timestamp 1681708930
transform 1 0 1036 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2817
timestamp 1681708930
transform 1 0 1044 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2843
timestamp 1681708930
transform 1 0 1012 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_2862
timestamp 1681708930
transform 1 0 1020 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2863
timestamp 1681708930
transform 1 0 1036 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2864
timestamp 1681708930
transform 1 0 1044 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2935
timestamp 1681708930
transform 1 0 1012 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2936
timestamp 1681708930
transform 1 0 1028 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2881
timestamp 1681708930
transform 1 0 1012 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2818
timestamp 1681708930
transform 1 0 1068 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2937
timestamp 1681708930
transform 1 0 1060 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2882
timestamp 1681708930
transform 1 0 1060 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_2981
timestamp 1681708930
transform 1 0 1068 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_2938
timestamp 1681708930
transform 1 0 1084 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2819
timestamp 1681708930
transform 1 0 1100 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_2775
timestamp 1681708930
transform 1 0 1140 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2819
timestamp 1681708930
transform 1 0 1140 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2820
timestamp 1681708930
transform 1 0 1172 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2865
timestamp 1681708930
transform 1 0 1108 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2866
timestamp 1681708930
transform 1 0 1124 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2867
timestamp 1681708930
transform 1 0 1140 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2939
timestamp 1681708930
transform 1 0 1124 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2883
timestamp 1681708930
transform 1 0 1124 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_2940
timestamp 1681708930
transform 1 0 1180 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2884
timestamp 1681708930
transform 1 0 1172 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2765
timestamp 1681708930
transform 1 0 1292 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2776
timestamp 1681708930
transform 1 0 1292 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2821
timestamp 1681708930
transform 1 0 1260 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2868
timestamp 1681708930
transform 1 0 1236 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2869
timestamp 1681708930
transform 1 0 1260 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2798
timestamp 1681708930
transform 1 0 1300 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_2941
timestamp 1681708930
transform 1 0 1292 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2822
timestamp 1681708930
transform 1 0 1340 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2942
timestamp 1681708930
transform 1 0 1340 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2943
timestamp 1681708930
transform 1 0 1348 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2885
timestamp 1681708930
transform 1 0 1348 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2900
timestamp 1681708930
transform 1 0 1300 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2901
timestamp 1681708930
transform 1 0 1316 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2777
timestamp 1681708930
transform 1 0 1412 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_2870
timestamp 1681708930
transform 1 0 1404 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2944
timestamp 1681708930
transform 1 0 1396 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2902
timestamp 1681708930
transform 1 0 1404 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2778
timestamp 1681708930
transform 1 0 1428 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_2871
timestamp 1681708930
transform 1 0 1420 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2945
timestamp 1681708930
transform 1 0 1428 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2886
timestamp 1681708930
transform 1 0 1420 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2823
timestamp 1681708930
transform 1 0 1476 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2820
timestamp 1681708930
transform 1 0 1484 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_2844
timestamp 1681708930
transform 1 0 1484 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_2946
timestamp 1681708930
transform 1 0 1484 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2807
timestamp 1681708930
transform 1 0 1508 0 1 835
box -2 -2 2 2
use M3_M2  M3_M2_2824
timestamp 1681708930
transform 1 0 1508 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2784
timestamp 1681708930
transform 1 0 1532 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_2808
timestamp 1681708930
transform 1 0 1572 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_2821
timestamp 1681708930
transform 1 0 1516 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_2825
timestamp 1681708930
transform 1 0 1540 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2826
timestamp 1681708930
transform 1 0 1556 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2822
timestamp 1681708930
transform 1 0 1564 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2823
timestamp 1681708930
transform 1 0 1588 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_2827
timestamp 1681708930
transform 1 0 1596 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2872
timestamp 1681708930
transform 1 0 1508 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2873
timestamp 1681708930
transform 1 0 1524 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2874
timestamp 1681708930
transform 1 0 1540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2875
timestamp 1681708930
transform 1 0 1556 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2868
timestamp 1681708930
transform 1 0 1508 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2845
timestamp 1681708930
transform 1 0 1564 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_2876
timestamp 1681708930
transform 1 0 1580 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2877
timestamp 1681708930
transform 1 0 1596 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2947
timestamp 1681708930
transform 1 0 1524 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2948
timestamp 1681708930
transform 1 0 1548 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2887
timestamp 1681708930
transform 1 0 1492 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2888
timestamp 1681708930
transform 1 0 1540 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2869
timestamp 1681708930
transform 1 0 1580 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_2878
timestamp 1681708930
transform 1 0 1612 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2846
timestamp 1681708930
transform 1 0 1620 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_2949
timestamp 1681708930
transform 1 0 1604 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2870
timestamp 1681708930
transform 1 0 1612 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2766
timestamp 1681708930
transform 1 0 1644 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2847
timestamp 1681708930
transform 1 0 1644 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_2950
timestamp 1681708930
transform 1 0 1636 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2951
timestamp 1681708930
transform 1 0 1644 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2828
timestamp 1681708930
transform 1 0 1660 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2982
timestamp 1681708930
transform 1 0 1660 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_2829
timestamp 1681708930
transform 1 0 1700 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2767
timestamp 1681708930
transform 1 0 1748 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2768
timestamp 1681708930
transform 1 0 1772 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2799
timestamp 1681708930
transform 1 0 1764 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2830
timestamp 1681708930
transform 1 0 1780 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2879
timestamp 1681708930
transform 1 0 1700 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2880
timestamp 1681708930
transform 1 0 1724 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2848
timestamp 1681708930
transform 1 0 1748 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_2881
timestamp 1681708930
transform 1 0 1756 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2952
timestamp 1681708930
transform 1 0 1716 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2889
timestamp 1681708930
transform 1 0 1724 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_2953
timestamp 1681708930
transform 1 0 1772 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2954
timestamp 1681708930
transform 1 0 1780 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2903
timestamp 1681708930
transform 1 0 1676 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2904
timestamp 1681708930
transform 1 0 1716 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2905
timestamp 1681708930
transform 1 0 1740 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2769
timestamp 1681708930
transform 1 0 1828 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2779
timestamp 1681708930
transform 1 0 1820 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2800
timestamp 1681708930
transform 1 0 1820 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2831
timestamp 1681708930
transform 1 0 1812 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2882
timestamp 1681708930
transform 1 0 1788 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2883
timestamp 1681708930
transform 1 0 1796 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2849
timestamp 1681708930
transform 1 0 1804 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2801
timestamp 1681708930
transform 1 0 1860 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_2884
timestamp 1681708930
transform 1 0 1812 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2885
timestamp 1681708930
transform 1 0 1828 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2886
timestamp 1681708930
transform 1 0 1836 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2887
timestamp 1681708930
transform 1 0 1852 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2871
timestamp 1681708930
transform 1 0 1796 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2850
timestamp 1681708930
transform 1 0 1860 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2785
timestamp 1681708930
transform 1 0 1876 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_2888
timestamp 1681708930
transform 1 0 1868 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2889
timestamp 1681708930
transform 1 0 1876 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2955
timestamp 1681708930
transform 1 0 1804 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2956
timestamp 1681708930
transform 1 0 1820 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2957
timestamp 1681708930
transform 1 0 1828 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2958
timestamp 1681708930
transform 1 0 1844 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2959
timestamp 1681708930
transform 1 0 1860 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2960
timestamp 1681708930
transform 1 0 1868 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2890
timestamp 1681708930
transform 1 0 1844 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2891
timestamp 1681708930
transform 1 0 1868 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2906
timestamp 1681708930
transform 1 0 1868 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2851
timestamp 1681708930
transform 1 0 1900 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_2890
timestamp 1681708930
transform 1 0 1932 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2852
timestamp 1681708930
transform 1 0 1940 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2770
timestamp 1681708930
transform 1 0 1964 0 1 865
box -3 -3 3 3
use M2_M1  M2_M1_2891
timestamp 1681708930
transform 1 0 1948 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2892
timestamp 1681708930
transform 1 0 1956 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2961
timestamp 1681708930
transform 1 0 1916 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2962
timestamp 1681708930
transform 1 0 1940 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2963
timestamp 1681708930
transform 1 0 1948 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2892
timestamp 1681708930
transform 1 0 1916 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2893
timestamp 1681708930
transform 1 0 1948 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2832
timestamp 1681708930
transform 1 0 2020 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2893
timestamp 1681708930
transform 1 0 1996 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2853
timestamp 1681708930
transform 1 0 2004 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_2894
timestamp 1681708930
transform 1 0 2020 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2895
timestamp 1681708930
transform 1 0 2028 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2964
timestamp 1681708930
transform 1 0 2004 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2965
timestamp 1681708930
transform 1 0 2012 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2966
timestamp 1681708930
transform 1 0 2036 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2907
timestamp 1681708930
transform 1 0 2036 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2833
timestamp 1681708930
transform 1 0 2068 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2896
timestamp 1681708930
transform 1 0 2068 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2897
timestamp 1681708930
transform 1 0 2092 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2854
timestamp 1681708930
transform 1 0 2100 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_2898
timestamp 1681708930
transform 1 0 2108 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2872
timestamp 1681708930
transform 1 0 2092 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2834
timestamp 1681708930
transform 1 0 2124 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2899
timestamp 1681708930
transform 1 0 2116 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2900
timestamp 1681708930
transform 1 0 2124 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2855
timestamp 1681708930
transform 1 0 2132 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2835
timestamp 1681708930
transform 1 0 2164 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2901
timestamp 1681708930
transform 1 0 2140 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2902
timestamp 1681708930
transform 1 0 2156 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2967
timestamp 1681708930
transform 1 0 2132 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2908
timestamp 1681708930
transform 1 0 2132 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_2968
timestamp 1681708930
transform 1 0 2196 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2809
timestamp 1681708930
transform 1 0 2228 0 1 835
box -2 -2 2 2
use M3_M2  M3_M2_2836
timestamp 1681708930
transform 1 0 2220 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2903
timestamp 1681708930
transform 1 0 2220 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2786
timestamp 1681708930
transform 1 0 2244 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2802
timestamp 1681708930
transform 1 0 2252 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_2824
timestamp 1681708930
transform 1 0 2236 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2825
timestamp 1681708930
transform 1 0 2244 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2969
timestamp 1681708930
transform 1 0 2228 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2837
timestamp 1681708930
transform 1 0 2260 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2904
timestamp 1681708930
transform 1 0 2244 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2970
timestamp 1681708930
transform 1 0 2244 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2909
timestamp 1681708930
transform 1 0 2244 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_2905
timestamp 1681708930
transform 1 0 2268 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2803
timestamp 1681708930
transform 1 0 2276 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_2826
timestamp 1681708930
transform 1 0 2276 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_2856
timestamp 1681708930
transform 1 0 2276 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2787
timestamp 1681708930
transform 1 0 2292 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_2827
timestamp 1681708930
transform 1 0 2316 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2906
timestamp 1681708930
transform 1 0 2308 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2971
timestamp 1681708930
transform 1 0 2292 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2873
timestamp 1681708930
transform 1 0 2300 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2857
timestamp 1681708930
transform 1 0 2316 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_2828
timestamp 1681708930
transform 1 0 2364 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2907
timestamp 1681708930
transform 1 0 2348 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2858
timestamp 1681708930
transform 1 0 2364 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_2908
timestamp 1681708930
transform 1 0 2380 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2972
timestamp 1681708930
transform 1 0 2356 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2973
timestamp 1681708930
transform 1 0 2364 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2974
timestamp 1681708930
transform 1 0 2396 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2829
timestamp 1681708930
transform 1 0 2412 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2975
timestamp 1681708930
transform 1 0 2428 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2771
timestamp 1681708930
transform 1 0 2436 0 1 865
box -3 -3 3 3
use M2_M1  M2_M1_2830
timestamp 1681708930
transform 1 0 2436 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2909
timestamp 1681708930
transform 1 0 2452 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_2838
timestamp 1681708930
transform 1 0 2476 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_2831
timestamp 1681708930
transform 1 0 2484 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2976
timestamp 1681708930
transform 1 0 2468 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2977
timestamp 1681708930
transform 1 0 2508 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2772
timestamp 1681708930
transform 1 0 2532 0 1 865
box -3 -3 3 3
use M2_M1  M2_M1_2978
timestamp 1681708930
transform 1 0 2540 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2894
timestamp 1681708930
transform 1 0 2548 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_2910
timestamp 1681708930
transform 1 0 2564 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2832
timestamp 1681708930
transform 1 0 2580 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_2839
timestamp 1681708930
transform 1 0 2596 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2859
timestamp 1681708930
transform 1 0 2580 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_2911
timestamp 1681708930
transform 1 0 2588 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2912
timestamp 1681708930
transform 1 0 2596 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2913
timestamp 1681708930
transform 1 0 2604 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2979
timestamp 1681708930
transform 1 0 2588 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2895
timestamp 1681708930
transform 1 0 2588 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2860
timestamp 1681708930
transform 1 0 2612 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_2914
timestamp 1681708930
transform 1 0 2660 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2980
timestamp 1681708930
transform 1 0 2612 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_2896
timestamp 1681708930
transform 1 0 2612 0 1 795
box -3 -3 3 3
use top_mod_new_VIA0  top_mod_new_VIA0_36
timestamp 1681708930
transform 1 0 48 0 1 770
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_69
timestamp 1681708930
transform -1 0 168 0 1 770
box -8 -3 104 105
use NAND2X1  NAND2X1_63
timestamp 1681708930
transform 1 0 168 0 1 770
box -8 -3 32 105
use OAI21X1  OAI21X1_68
timestamp 1681708930
transform -1 0 224 0 1 770
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_71
timestamp 1681708930
transform 1 0 224 0 1 770
box -8 -3 104 105
use FILL  FILL_1133
timestamp 1681708930
transform 1 0 320 0 1 770
box -8 -3 16 105
use AND2X2  AND2X2_4
timestamp 1681708930
transform -1 0 360 0 1 770
box -8 -3 40 105
use INVX2  INVX2_181
timestamp 1681708930
transform -1 0 376 0 1 770
box -9 -3 26 105
use INVX2  INVX2_182
timestamp 1681708930
transform -1 0 392 0 1 770
box -9 -3 26 105
use INVX2  INVX2_183
timestamp 1681708930
transform 1 0 392 0 1 770
box -9 -3 26 105
use FILL  FILL_1134
timestamp 1681708930
transform 1 0 408 0 1 770
box -8 -3 16 105
use INVX2  INVX2_184
timestamp 1681708930
transform -1 0 432 0 1 770
box -9 -3 26 105
use INVX2  INVX2_185
timestamp 1681708930
transform 1 0 432 0 1 770
box -9 -3 26 105
use FILL  FILL_1135
timestamp 1681708930
transform 1 0 448 0 1 770
box -8 -3 16 105
use FILL  FILL_1154
timestamp 1681708930
transform 1 0 456 0 1 770
box -8 -3 16 105
use FILL  FILL_1155
timestamp 1681708930
transform 1 0 464 0 1 770
box -8 -3 16 105
use FILL  FILL_1156
timestamp 1681708930
transform 1 0 472 0 1 770
box -8 -3 16 105
use FILL  FILL_1157
timestamp 1681708930
transform 1 0 480 0 1 770
box -8 -3 16 105
use INVX2  INVX2_188
timestamp 1681708930
transform -1 0 504 0 1 770
box -9 -3 26 105
use NAND2X1  NAND2X1_66
timestamp 1681708930
transform 1 0 504 0 1 770
box -8 -3 32 105
use FILL  FILL_1158
timestamp 1681708930
transform 1 0 528 0 1 770
box -8 -3 16 105
use FILL  FILL_1159
timestamp 1681708930
transform 1 0 536 0 1 770
box -8 -3 16 105
use FILL  FILL_1160
timestamp 1681708930
transform 1 0 544 0 1 770
box -8 -3 16 105
use FILL  FILL_1161
timestamp 1681708930
transform 1 0 552 0 1 770
box -8 -3 16 105
use FILL  FILL_1162
timestamp 1681708930
transform 1 0 560 0 1 770
box -8 -3 16 105
use FILL  FILL_1163
timestamp 1681708930
transform 1 0 568 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_64
timestamp 1681708930
transform 1 0 576 0 1 770
box -8 -3 46 105
use FILL  FILL_1164
timestamp 1681708930
transform 1 0 616 0 1 770
box -8 -3 16 105
use FILL  FILL_1167
timestamp 1681708930
transform 1 0 624 0 1 770
box -8 -3 16 105
use FILL  FILL_1168
timestamp 1681708930
transform 1 0 632 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_2910
timestamp 1681708930
transform 1 0 652 0 1 775
box -3 -3 3 3
use FILL  FILL_1169
timestamp 1681708930
transform 1 0 640 0 1 770
box -8 -3 16 105
use INVX2  INVX2_189
timestamp 1681708930
transform 1 0 648 0 1 770
box -9 -3 26 105
use FILL  FILL_1170
timestamp 1681708930
transform 1 0 664 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_2911
timestamp 1681708930
transform 1 0 684 0 1 775
box -3 -3 3 3
use NAND3X1  NAND3X1_107
timestamp 1681708930
transform 1 0 672 0 1 770
box -8 -3 40 105
use AOI22X1  AOI22X1_66
timestamp 1681708930
transform -1 0 744 0 1 770
box -8 -3 46 105
use FILL  FILL_1173
timestamp 1681708930
transform 1 0 744 0 1 770
box -8 -3 16 105
use FILL  FILL_1177
timestamp 1681708930
transform 1 0 752 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_2912
timestamp 1681708930
transform 1 0 796 0 1 775
box -3 -3 3 3
use XOR2X1  XOR2X1_152
timestamp 1681708930
transform -1 0 816 0 1 770
box -8 -3 64 105
use M3_M2  M3_M2_2913
timestamp 1681708930
transform 1 0 828 0 1 775
box -3 -3 3 3
use OAI21X1  OAI21X1_71
timestamp 1681708930
transform -1 0 848 0 1 770
box -8 -3 34 105
use FILL  FILL_1178
timestamp 1681708930
transform 1 0 848 0 1 770
box -8 -3 16 105
use FILL  FILL_1189
timestamp 1681708930
transform 1 0 856 0 1 770
box -8 -3 16 105
use INVX2  INVX2_192
timestamp 1681708930
transform 1 0 864 0 1 770
box -9 -3 26 105
use FILL  FILL_1191
timestamp 1681708930
transform 1 0 880 0 1 770
box -8 -3 16 105
use FILL  FILL_1192
timestamp 1681708930
transform 1 0 888 0 1 770
box -8 -3 16 105
use FILL  FILL_1193
timestamp 1681708930
transform 1 0 896 0 1 770
box -8 -3 16 105
use FILL  FILL_1194
timestamp 1681708930
transform 1 0 904 0 1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_108
timestamp 1681708930
transform 1 0 912 0 1 770
box -8 -3 40 105
use FILL  FILL_1195
timestamp 1681708930
transform 1 0 944 0 1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_109
timestamp 1681708930
transform -1 0 984 0 1 770
box -8 -3 40 105
use FILL  FILL_1196
timestamp 1681708930
transform 1 0 984 0 1 770
box -8 -3 16 105
use FILL  FILL_1202
timestamp 1681708930
transform 1 0 992 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_68
timestamp 1681708930
transform -1 0 1040 0 1 770
box -8 -3 46 105
use OR2X1  OR2X1_19
timestamp 1681708930
transform -1 0 1072 0 1 770
box -8 -3 40 105
use FILL  FILL_1203
timestamp 1681708930
transform 1 0 1072 0 1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_69
timestamp 1681708930
transform 1 0 1080 0 1 770
box -8 -3 32 105
use M3_M2  M3_M2_2914
timestamp 1681708930
transform 1 0 1132 0 1 775
box -3 -3 3 3
use INVX2  INVX2_194
timestamp 1681708930
transform 1 0 1104 0 1 770
box -9 -3 26 105
use M3_M2  M3_M2_2915
timestamp 1681708930
transform 1 0 1180 0 1 775
box -3 -3 3 3
use XNOR2X1  XNOR2X1_47
timestamp 1681708930
transform -1 0 1176 0 1 770
box -8 -3 64 105
use M3_M2  M3_M2_2916
timestamp 1681708930
transform 1 0 1228 0 1 775
box -3 -3 3 3
use XOR2X1  XOR2X1_153
timestamp 1681708930
transform -1 0 1232 0 1 770
box -8 -3 64 105
use XOR2X1  XOR2X1_154
timestamp 1681708930
transform 1 0 1232 0 1 770
box -8 -3 64 105
use XOR2X1  XOR2X1_155
timestamp 1681708930
transform -1 0 1344 0 1 770
box -8 -3 64 105
use XOR2X1  XOR2X1_156
timestamp 1681708930
transform 1 0 1344 0 1 770
box -8 -3 64 105
use FILL  FILL_1211
timestamp 1681708930
transform 1 0 1400 0 1 770
box -8 -3 16 105
use FILL  FILL_1212
timestamp 1681708930
transform 1 0 1408 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_2917
timestamp 1681708930
transform 1 0 1428 0 1 775
box -3 -3 3 3
use FILL  FILL_1213
timestamp 1681708930
transform 1 0 1416 0 1 770
box -8 -3 16 105
use XOR2X1  XOR2X1_157
timestamp 1681708930
transform -1 0 1480 0 1 770
box -8 -3 64 105
use FILL  FILL_1214
timestamp 1681708930
transform 1 0 1480 0 1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_112
timestamp 1681708930
transform -1 0 1520 0 1 770
box -8 -3 40 105
use AOI22X1  AOI22X1_69
timestamp 1681708930
transform 1 0 1520 0 1 770
box -8 -3 46 105
use NAND3X1  NAND3X1_113
timestamp 1681708930
transform -1 0 1592 0 1 770
box -8 -3 40 105
use INVX2  INVX2_195
timestamp 1681708930
transform -1 0 1608 0 1 770
box -9 -3 26 105
use FILL  FILL_1215
timestamp 1681708930
transform 1 0 1608 0 1 770
box -8 -3 16 105
use OR2X1  OR2X1_20
timestamp 1681708930
transform -1 0 1648 0 1 770
box -8 -3 40 105
use FILL  FILL_1216
timestamp 1681708930
transform 1 0 1648 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_2918
timestamp 1681708930
transform 1 0 1668 0 1 775
box -3 -3 3 3
use FILL  FILL_1233
timestamp 1681708930
transform 1 0 1656 0 1 770
box -8 -3 16 105
use XNOR2X1  XNOR2X1_48
timestamp 1681708930
transform 1 0 1664 0 1 770
box -8 -3 64 105
use M3_M2  M3_M2_2919
timestamp 1681708930
transform 1 0 1772 0 1 775
box -3 -3 3 3
use XOR2X1  XOR2X1_164
timestamp 1681708930
transform 1 0 1720 0 1 770
box -8 -3 64 105
use INVX2  INVX2_198
timestamp 1681708930
transform 1 0 1776 0 1 770
box -9 -3 26 105
use AOI22X1  AOI22X1_71
timestamp 1681708930
transform -1 0 1832 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_72
timestamp 1681708930
transform -1 0 1872 0 1 770
box -8 -3 46 105
use FILL  FILL_1234
timestamp 1681708930
transform 1 0 1872 0 1 770
box -8 -3 16 105
use FILL  FILL_1235
timestamp 1681708930
transform 1 0 1880 0 1 770
box -8 -3 16 105
use FILL  FILL_1236
timestamp 1681708930
transform 1 0 1888 0 1 770
box -8 -3 16 105
use FILL  FILL_1237
timestamp 1681708930
transform 1 0 1896 0 1 770
box -8 -3 16 105
use FILL  FILL_1238
timestamp 1681708930
transform 1 0 1904 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_73
timestamp 1681708930
transform -1 0 1952 0 1 770
box -8 -3 46 105
use FILL  FILL_1239
timestamp 1681708930
transform 1 0 1952 0 1 770
box -8 -3 16 105
use FILL  FILL_1240
timestamp 1681708930
transform 1 0 1960 0 1 770
box -8 -3 16 105
use FILL  FILL_1241
timestamp 1681708930
transform 1 0 1968 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_74
timestamp 1681708930
transform -1 0 2016 0 1 770
box -8 -3 46 105
use INVX2  INVX2_199
timestamp 1681708930
transform 1 0 2016 0 1 770
box -9 -3 26 105
use FILL  FILL_1242
timestamp 1681708930
transform 1 0 2032 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_2920
timestamp 1681708930
transform 1 0 2060 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2921
timestamp 1681708930
transform 1 0 2100 0 1 775
box -3 -3 3 3
use XOR2X1  XOR2X1_165
timestamp 1681708930
transform 1 0 2040 0 1 770
box -8 -3 64 105
use FILL  FILL_1243
timestamp 1681708930
transform 1 0 2096 0 1 770
box -8 -3 16 105
use INVX2  INVX2_200
timestamp 1681708930
transform 1 0 2104 0 1 770
box -9 -3 26 105
use AOI22X1  AOI22X1_75
timestamp 1681708930
transform -1 0 2160 0 1 770
box -8 -3 46 105
use FILL  FILL_1244
timestamp 1681708930
transform 1 0 2160 0 1 770
box -8 -3 16 105
use FILL  FILL_1245
timestamp 1681708930
transform 1 0 2168 0 1 770
box -8 -3 16 105
use FILL  FILL_1250
timestamp 1681708930
transform 1 0 2176 0 1 770
box -8 -3 16 105
use INVX2  INVX2_204
timestamp 1681708930
transform -1 0 2200 0 1 770
box -9 -3 26 105
use NOR2X1  NOR2X1_65
timestamp 1681708930
transform 1 0 2200 0 1 770
box -8 -3 32 105
use FILL  FILL_1251
timestamp 1681708930
transform 1 0 2224 0 1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_116
timestamp 1681708930
transform 1 0 2232 0 1 770
box -8 -3 40 105
use FILL  FILL_1255
timestamp 1681708930
transform 1 0 2264 0 1 770
box -8 -3 16 105
use FILL  FILL_1256
timestamp 1681708930
transform 1 0 2272 0 1 770
box -8 -3 16 105
use AOI21X1  AOI21X1_40
timestamp 1681708930
transform 1 0 2280 0 1 770
box -7 -3 39 105
use FILL  FILL_1257
timestamp 1681708930
transform 1 0 2312 0 1 770
box -8 -3 16 105
use FILL  FILL_1258
timestamp 1681708930
transform 1 0 2320 0 1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_72
timestamp 1681708930
transform -1 0 2360 0 1 770
box -8 -3 34 105
use M3_M2  M3_M2_2922
timestamp 1681708930
transform 1 0 2396 0 1 775
box -3 -3 3 3
use OAI21X1  OAI21X1_73
timestamp 1681708930
transform -1 0 2392 0 1 770
box -8 -3 34 105
use NAND2X1  NAND2X1_70
timestamp 1681708930
transform 1 0 2392 0 1 770
box -8 -3 32 105
use FILL  FILL_1259
timestamp 1681708930
transform 1 0 2416 0 1 770
box -8 -3 16 105
use FILL  FILL_1260
timestamp 1681708930
transform 1 0 2424 0 1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_74
timestamp 1681708930
transform -1 0 2464 0 1 770
box -8 -3 34 105
use NAND2X1  NAND2X1_71
timestamp 1681708930
transform 1 0 2464 0 1 770
box -8 -3 32 105
use FILL  FILL_1261
timestamp 1681708930
transform 1 0 2488 0 1 770
box -8 -3 16 105
use FILL  FILL_1262
timestamp 1681708930
transform 1 0 2496 0 1 770
box -8 -3 16 105
use FILL  FILL_1263
timestamp 1681708930
transform 1 0 2504 0 1 770
box -8 -3 16 105
use INVX2  INVX2_205
timestamp 1681708930
transform 1 0 2512 0 1 770
box -9 -3 26 105
use FILL  FILL_1264
timestamp 1681708930
transform 1 0 2528 0 1 770
box -8 -3 16 105
use FILL  FILL_1265
timestamp 1681708930
transform 1 0 2536 0 1 770
box -8 -3 16 105
use FILL  FILL_1266
timestamp 1681708930
transform 1 0 2544 0 1 770
box -8 -3 16 105
use FILL  FILL_1267
timestamp 1681708930
transform 1 0 2552 0 1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_72
timestamp 1681708930
transform 1 0 2560 0 1 770
box -8 -3 32 105
use INVX2  INVX2_206
timestamp 1681708930
transform 1 0 2584 0 1 770
box -9 -3 26 105
use FILL  FILL_1268
timestamp 1681708930
transform 1 0 2600 0 1 770
box -8 -3 16 105
use XOR2X1  XOR2X1_166
timestamp 1681708930
transform -1 0 2664 0 1 770
box -8 -3 64 105
use top_mod_new_VIA0  top_mod_new_VIA0_37
timestamp 1681708930
transform 1 0 2688 0 1 770
box -10 -3 10 3
use M3_M2  M3_M2_2956
timestamp 1681708930
transform 1 0 132 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2937
timestamp 1681708930
transform 1 0 196 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2957
timestamp 1681708930
transform 1 0 188 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_2984
timestamp 1681708930
transform 1 0 156 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2985
timestamp 1681708930
transform 1 0 172 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2986
timestamp 1681708930
transform 1 0 188 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3047
timestamp 1681708930
transform 1 0 76 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3048
timestamp 1681708930
transform 1 0 132 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3013
timestamp 1681708930
transform 1 0 76 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3014
timestamp 1681708930
transform 1 0 172 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2978
timestamp 1681708930
transform 1 0 196 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2979
timestamp 1681708930
transform 1 0 212 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_2987
timestamp 1681708930
transform 1 0 220 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3108
timestamp 1681708930
transform 1 0 188 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2988
timestamp 1681708930
transform 1 0 260 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_2980
timestamp 1681708930
transform 1 0 276 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_3049
timestamp 1681708930
transform 1 0 268 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3050
timestamp 1681708930
transform 1 0 276 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3033
timestamp 1681708930
transform 1 0 300 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2923
timestamp 1681708930
transform 1 0 324 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_2989
timestamp 1681708930
transform 1 0 316 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_2981
timestamp 1681708930
transform 1 0 332 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_2990
timestamp 1681708930
transform 1 0 348 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3051
timestamp 1681708930
transform 1 0 332 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2991
timestamp 1681708930
transform 1 0 356 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3034
timestamp 1681708930
transform 1 0 356 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2982
timestamp 1681708930
transform 1 0 380 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_3109
timestamp 1681708930
transform 1 0 380 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3035
timestamp 1681708930
transform 1 0 380 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2924
timestamp 1681708930
transform 1 0 404 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_3052
timestamp 1681708930
transform 1 0 396 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3110
timestamp 1681708930
transform 1 0 404 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3054
timestamp 1681708930
transform 1 0 404 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_2992
timestamp 1681708930
transform 1 0 444 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_2938
timestamp 1681708930
transform 1 0 516 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_2993
timestamp 1681708930
transform 1 0 468 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2994
timestamp 1681708930
transform 1 0 484 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_2983
timestamp 1681708930
transform 1 0 492 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2984
timestamp 1681708930
transform 1 0 508 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_2995
timestamp 1681708930
transform 1 0 516 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2996
timestamp 1681708930
transform 1 0 524 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3053
timestamp 1681708930
transform 1 0 460 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3054
timestamp 1681708930
transform 1 0 476 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_2996
timestamp 1681708930
transform 1 0 484 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_3055
timestamp 1681708930
transform 1 0 492 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_2997
timestamp 1681708930
transform 1 0 500 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_3111
timestamp 1681708930
transform 1 0 500 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3036
timestamp 1681708930
transform 1 0 476 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3055
timestamp 1681708930
transform 1 0 500 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3066
timestamp 1681708930
transform 1 0 468 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3067
timestamp 1681708930
transform 1 0 484 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_3056
timestamp 1681708930
transform 1 0 540 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3057
timestamp 1681708930
transform 1 0 548 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3037
timestamp 1681708930
transform 1 0 540 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_2997
timestamp 1681708930
transform 1 0 604 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3112
timestamp 1681708930
transform 1 0 620 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3128
timestamp 1681708930
transform 1 0 596 0 1 705
box -2 -2 2 2
use M3_M2  M3_M2_3038
timestamp 1681708930
transform 1 0 612 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_3058
timestamp 1681708930
transform 1 0 636 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2998
timestamp 1681708930
transform 1 0 644 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3059
timestamp 1681708930
transform 1 0 644 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2999
timestamp 1681708930
transform 1 0 676 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3000
timestamp 1681708930
transform 1 0 692 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3060
timestamp 1681708930
transform 1 0 716 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3001
timestamp 1681708930
transform 1 0 748 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_2985
timestamp 1681708930
transform 1 0 772 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_3056
timestamp 1681708930
transform 1 0 812 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2925
timestamp 1681708930
transform 1 0 836 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_3113
timestamp 1681708930
transform 1 0 828 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3002
timestamp 1681708930
transform 1 0 852 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3039
timestamp 1681708930
transform 1 0 844 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_3061
timestamp 1681708930
transform 1 0 868 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3015
timestamp 1681708930
transform 1 0 868 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2939
timestamp 1681708930
transform 1 0 900 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2940
timestamp 1681708930
transform 1 0 916 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2958
timestamp 1681708930
transform 1 0 884 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_3062
timestamp 1681708930
transform 1 0 884 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3114
timestamp 1681708930
transform 1 0 876 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3040
timestamp 1681708930
transform 1 0 860 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_3063
timestamp 1681708930
transform 1 0 916 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3064
timestamp 1681708930
transform 1 0 924 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3115
timestamp 1681708930
transform 1 0 908 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3016
timestamp 1681708930
transform 1 0 916 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3041
timestamp 1681708930
transform 1 0 924 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2941
timestamp 1681708930
transform 1 0 956 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2959
timestamp 1681708930
transform 1 0 972 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_3003
timestamp 1681708930
transform 1 0 956 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3004
timestamp 1681708930
transform 1 0 972 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_2998
timestamp 1681708930
transform 1 0 948 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_3065
timestamp 1681708930
transform 1 0 964 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3057
timestamp 1681708930
transform 1 0 940 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3017
timestamp 1681708930
transform 1 0 964 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_3066
timestamp 1681708930
transform 1 0 988 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3116
timestamp 1681708930
transform 1 0 988 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_2926
timestamp 1681708930
transform 1 0 1020 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2927
timestamp 1681708930
transform 1 0 1044 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_3005
timestamp 1681708930
transform 1 0 1044 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_2999
timestamp 1681708930
transform 1 0 1028 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_3117
timestamp 1681708930
transform 1 0 1044 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3129
timestamp 1681708930
transform 1 0 1036 0 1 705
box -2 -2 2 2
use M3_M2  M3_M2_3042
timestamp 1681708930
transform 1 0 1044 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3058
timestamp 1681708930
transform 1 0 1036 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2928
timestamp 1681708930
transform 1 0 1068 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2960
timestamp 1681708930
transform 1 0 1060 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_3067
timestamp 1681708930
transform 1 0 1060 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_2942
timestamp 1681708930
transform 1 0 1084 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_3006
timestamp 1681708930
transform 1 0 1108 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3068
timestamp 1681708930
transform 1 0 1100 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3059
timestamp 1681708930
transform 1 0 1108 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_3007
timestamp 1681708930
transform 1 0 1124 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_2943
timestamp 1681708930
transform 1 0 1140 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2944
timestamp 1681708930
transform 1 0 1172 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2945
timestamp 1681708930
transform 1 0 1204 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_3008
timestamp 1681708930
transform 1 0 1148 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3069
timestamp 1681708930
transform 1 0 1140 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_2961
timestamp 1681708930
transform 1 0 1196 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_3009
timestamp 1681708930
transform 1 0 1196 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3010
timestamp 1681708930
transform 1 0 1204 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_2929
timestamp 1681708930
transform 1 0 1252 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2946
timestamp 1681708930
transform 1 0 1300 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2962
timestamp 1681708930
transform 1 0 1260 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_3011
timestamp 1681708930
transform 1 0 1252 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3012
timestamp 1681708930
transform 1 0 1260 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3070
timestamp 1681708930
transform 1 0 1228 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_2930
timestamp 1681708930
transform 1 0 1348 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_3013
timestamp 1681708930
transform 1 0 1308 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3014
timestamp 1681708930
transform 1 0 1316 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3071
timestamp 1681708930
transform 1 0 1284 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_2947
timestamp 1681708930
transform 1 0 1364 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_3015
timestamp 1681708930
transform 1 0 1372 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3072
timestamp 1681708930
transform 1 0 1340 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3018
timestamp 1681708930
transform 1 0 1316 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3043
timestamp 1681708930
transform 1 0 1300 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3000
timestamp 1681708930
transform 1 0 1364 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_3016
timestamp 1681708930
transform 1 0 1420 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3017
timestamp 1681708930
transform 1 0 1428 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3073
timestamp 1681708930
transform 1 0 1396 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3074
timestamp 1681708930
transform 1 0 1404 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3019
timestamp 1681708930
transform 1 0 1372 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3020
timestamp 1681708930
transform 1 0 1404 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3044
timestamp 1681708930
transform 1 0 1396 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_3075
timestamp 1681708930
transform 1 0 1476 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_2963
timestamp 1681708930
transform 1 0 1492 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_3018
timestamp 1681708930
transform 1 0 1492 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_2948
timestamp 1681708930
transform 1 0 1516 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2949
timestamp 1681708930
transform 1 0 1548 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2964
timestamp 1681708930
transform 1 0 1516 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2965
timestamp 1681708930
transform 1 0 1540 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_3019
timestamp 1681708930
transform 1 0 1516 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3020
timestamp 1681708930
transform 1 0 1532 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3021
timestamp 1681708930
transform 1 0 1540 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3076
timestamp 1681708930
transform 1 0 1508 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3077
timestamp 1681708930
transform 1 0 1524 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3078
timestamp 1681708930
transform 1 0 1540 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3021
timestamp 1681708930
transform 1 0 1508 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3022
timestamp 1681708930
transform 1 0 1540 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3045
timestamp 1681708930
transform 1 0 1516 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3068
timestamp 1681708930
transform 1 0 1532 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2966
timestamp 1681708930
transform 1 0 1564 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_3022
timestamp 1681708930
transform 1 0 1556 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3023
timestamp 1681708930
transform 1 0 1572 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3024
timestamp 1681708930
transform 1 0 1588 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3079
timestamp 1681708930
transform 1 0 1564 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3080
timestamp 1681708930
transform 1 0 1580 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3023
timestamp 1681708930
transform 1 0 1556 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3046
timestamp 1681708930
transform 1 0 1548 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3047
timestamp 1681708930
transform 1 0 1564 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2931
timestamp 1681708930
transform 1 0 1604 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_3081
timestamp 1681708930
transform 1 0 1604 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3118
timestamp 1681708930
transform 1 0 1612 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3048
timestamp 1681708930
transform 1 0 1612 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3069
timestamp 1681708930
transform 1 0 1652 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2932
timestamp 1681708930
transform 1 0 1684 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_3082
timestamp 1681708930
transform 1 0 1668 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_2986
timestamp 1681708930
transform 1 0 1692 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_3083
timestamp 1681708930
transform 1 0 1692 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3119
timestamp 1681708930
transform 1 0 1684 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3130
timestamp 1681708930
transform 1 0 1676 0 1 705
box -2 -2 2 2
use M3_M2  M3_M2_2933
timestamp 1681708930
transform 1 0 1852 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2934
timestamp 1681708930
transform 1 0 1876 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2935
timestamp 1681708930
transform 1 0 1924 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2967
timestamp 1681708930
transform 1 0 1732 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2968
timestamp 1681708930
transform 1 0 1820 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_3025
timestamp 1681708930
transform 1 0 1732 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_2987
timestamp 1681708930
transform 1 0 1780 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_3026
timestamp 1681708930
transform 1 0 1820 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_2988
timestamp 1681708930
transform 1 0 1836 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2969
timestamp 1681708930
transform 1 0 1860 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2970
timestamp 1681708930
transform 1 0 1932 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_3027
timestamp 1681708930
transform 1 0 1844 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3028
timestamp 1681708930
transform 1 0 1932 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3029
timestamp 1681708930
transform 1 0 1948 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3084
timestamp 1681708930
transform 1 0 1740 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3085
timestamp 1681708930
transform 1 0 1788 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3086
timestamp 1681708930
transform 1 0 1836 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3087
timestamp 1681708930
transform 1 0 1844 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3088
timestamp 1681708930
transform 1 0 1852 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3001
timestamp 1681708930
transform 1 0 1868 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2936
timestamp 1681708930
transform 1 0 1996 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2971
timestamp 1681708930
transform 1 0 2044 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_3030
timestamp 1681708930
transform 1 0 2044 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3089
timestamp 1681708930
transform 1 0 1908 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3090
timestamp 1681708930
transform 1 0 1948 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3091
timestamp 1681708930
transform 1 0 1964 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3092
timestamp 1681708930
transform 1 0 2020 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3024
timestamp 1681708930
transform 1 0 1908 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3025
timestamp 1681708930
transform 1 0 1948 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3002
timestamp 1681708930
transform 1 0 2044 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2950
timestamp 1681708930
transform 1 0 2108 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2951
timestamp 1681708930
transform 1 0 2148 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2952
timestamp 1681708930
transform 1 0 2164 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2972
timestamp 1681708930
transform 1 0 2140 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_3031
timestamp 1681708930
transform 1 0 2140 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_2973
timestamp 1681708930
transform 1 0 2172 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_3032
timestamp 1681708930
transform 1 0 2164 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3093
timestamp 1681708930
transform 1 0 2060 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3049
timestamp 1681708930
transform 1 0 1996 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3003
timestamp 1681708930
transform 1 0 2108 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_3094
timestamp 1681708930
transform 1 0 2116 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3004
timestamp 1681708930
transform 1 0 2140 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_3095
timestamp 1681708930
transform 1 0 2156 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3096
timestamp 1681708930
transform 1 0 2164 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3050
timestamp 1681708930
transform 1 0 2148 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3070
timestamp 1681708930
transform 1 0 2084 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3060
timestamp 1681708930
transform 1 0 2164 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2953
timestamp 1681708930
transform 1 0 2188 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_3033
timestamp 1681708930
transform 1 0 2188 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3005
timestamp 1681708930
transform 1 0 2196 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_3120
timestamp 1681708930
transform 1 0 2204 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3131
timestamp 1681708930
transform 1 0 2196 0 1 705
box -2 -2 2 2
use M3_M2  M3_M2_3071
timestamp 1681708930
transform 1 0 2180 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2954
timestamp 1681708930
transform 1 0 2220 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2974
timestamp 1681708930
transform 1 0 2220 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_3121
timestamp 1681708930
transform 1 0 2220 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3132
timestamp 1681708930
transform 1 0 2212 0 1 705
box -2 -2 2 2
use M3_M2  M3_M2_3061
timestamp 1681708930
transform 1 0 2212 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2989
timestamp 1681708930
transform 1 0 2236 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_3034
timestamp 1681708930
transform 1 0 2268 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_2990
timestamp 1681708930
transform 1 0 2276 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_2983
timestamp 1681708930
transform 1 0 2292 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_3035
timestamp 1681708930
transform 1 0 2284 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3097
timestamp 1681708930
transform 1 0 2244 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3133
timestamp 1681708930
transform 1 0 2236 0 1 705
box -2 -2 2 2
use M3_M2  M3_M2_3006
timestamp 1681708930
transform 1 0 2260 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_3098
timestamp 1681708930
transform 1 0 2268 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3122
timestamp 1681708930
transform 1 0 2260 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3026
timestamp 1681708930
transform 1 0 2268 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_3099
timestamp 1681708930
transform 1 0 2284 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3051
timestamp 1681708930
transform 1 0 2284 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_3036
timestamp 1681708930
transform 1 0 2324 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_2975
timestamp 1681708930
transform 1 0 2348 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2991
timestamp 1681708930
transform 1 0 2340 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_3037
timestamp 1681708930
transform 1 0 2348 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3007
timestamp 1681708930
transform 1 0 2332 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_3100
timestamp 1681708930
transform 1 0 2340 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3101
timestamp 1681708930
transform 1 0 2356 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3027
timestamp 1681708930
transform 1 0 2324 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3062
timestamp 1681708930
transform 1 0 2316 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3028
timestamp 1681708930
transform 1 0 2340 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_3123
timestamp 1681708930
transform 1 0 2348 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3063
timestamp 1681708930
transform 1 0 2348 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3008
timestamp 1681708930
transform 1 0 2364 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_3124
timestamp 1681708930
transform 1 0 2364 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3052
timestamp 1681708930
transform 1 0 2364 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2992
timestamp 1681708930
transform 1 0 2380 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_3038
timestamp 1681708930
transform 1 0 2396 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3009
timestamp 1681708930
transform 1 0 2388 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3029
timestamp 1681708930
transform 1 0 2404 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2976
timestamp 1681708930
transform 1 0 2444 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_3039
timestamp 1681708930
transform 1 0 2420 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3053
timestamp 1681708930
transform 1 0 2412 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2993
timestamp 1681708930
transform 1 0 2428 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_3040
timestamp 1681708930
transform 1 0 2444 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3010
timestamp 1681708930
transform 1 0 2428 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_3041
timestamp 1681708930
transform 1 0 2492 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_2994
timestamp 1681708930
transform 1 0 2500 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_3102
timestamp 1681708930
transform 1 0 2436 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3103
timestamp 1681708930
transform 1 0 2468 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3011
timestamp 1681708930
transform 1 0 2500 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2955
timestamp 1681708930
transform 1 0 2540 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_3042
timestamp 1681708930
transform 1 0 2532 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3104
timestamp 1681708930
transform 1 0 2508 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3105
timestamp 1681708930
transform 1 0 2532 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3125
timestamp 1681708930
transform 1 0 2436 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3030
timestamp 1681708930
transform 1 0 2468 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_3126
timestamp 1681708930
transform 1 0 2508 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3127
timestamp 1681708930
transform 1 0 2524 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3134
timestamp 1681708930
transform 1 0 2516 0 1 705
box -2 -2 2 2
use M3_M2  M3_M2_3064
timestamp 1681708930
transform 1 0 2516 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2977
timestamp 1681708930
transform 1 0 2604 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_3043
timestamp 1681708930
transform 1 0 2580 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3044
timestamp 1681708930
transform 1 0 2588 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_2995
timestamp 1681708930
transform 1 0 2596 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_3045
timestamp 1681708930
transform 1 0 2604 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3106
timestamp 1681708930
transform 1 0 2604 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3107
timestamp 1681708930
transform 1 0 2620 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3031
timestamp 1681708930
transform 1 0 2588 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3065
timestamp 1681708930
transform 1 0 2588 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3012
timestamp 1681708930
transform 1 0 2628 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3032
timestamp 1681708930
transform 1 0 2620 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_3046
timestamp 1681708930
transform 1 0 2668 0 1 735
box -2 -2 2 2
use top_mod_new_VIA0  top_mod_new_VIA0_38
timestamp 1681708930
transform 1 0 24 0 1 670
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_70
timestamp 1681708930
transform -1 0 168 0 -1 770
box -8 -3 104 105
use NAND2X1  NAND2X1_64
timestamp 1681708930
transform 1 0 168 0 -1 770
box -8 -3 32 105
use OAI21X1  OAI21X1_69
timestamp 1681708930
transform -1 0 224 0 -1 770
box -8 -3 34 105
use INVX2  INVX2_186
timestamp 1681708930
transform -1 0 240 0 -1 770
box -9 -3 26 105
use FILL  FILL_1136
timestamp 1681708930
transform 1 0 240 0 -1 770
box -8 -3 16 105
use FILL  FILL_1137
timestamp 1681708930
transform 1 0 248 0 -1 770
box -8 -3 16 105
use FILL  FILL_1138
timestamp 1681708930
transform 1 0 256 0 -1 770
box -8 -3 16 105
use FILL  FILL_1139
timestamp 1681708930
transform 1 0 264 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_187
timestamp 1681708930
transform -1 0 288 0 -1 770
box -9 -3 26 105
use FILL  FILL_1140
timestamp 1681708930
transform 1 0 288 0 -1 770
box -8 -3 16 105
use FILL  FILL_1141
timestamp 1681708930
transform 1 0 296 0 -1 770
box -8 -3 16 105
use FILL  FILL_1142
timestamp 1681708930
transform 1 0 304 0 -1 770
box -8 -3 16 105
use FILL  FILL_1143
timestamp 1681708930
transform 1 0 312 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_70
timestamp 1681708930
transform 1 0 320 0 -1 770
box -8 -3 34 105
use FILL  FILL_1144
timestamp 1681708930
transform 1 0 352 0 -1 770
box -8 -3 16 105
use FILL  FILL_1145
timestamp 1681708930
transform 1 0 360 0 -1 770
box -8 -3 16 105
use FILL  FILL_1146
timestamp 1681708930
transform 1 0 368 0 -1 770
box -8 -3 16 105
use FILL  FILL_1147
timestamp 1681708930
transform 1 0 376 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_65
timestamp 1681708930
transform 1 0 384 0 -1 770
box -8 -3 32 105
use FILL  FILL_1148
timestamp 1681708930
transform 1 0 408 0 -1 770
box -8 -3 16 105
use FILL  FILL_1149
timestamp 1681708930
transform 1 0 416 0 -1 770
box -8 -3 16 105
use FILL  FILL_1150
timestamp 1681708930
transform 1 0 424 0 -1 770
box -8 -3 16 105
use FILL  FILL_1151
timestamp 1681708930
transform 1 0 432 0 -1 770
box -8 -3 16 105
use FILL  FILL_1152
timestamp 1681708930
transform 1 0 440 0 -1 770
box -8 -3 16 105
use FILL  FILL_1153
timestamp 1681708930
transform 1 0 448 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_65
timestamp 1681708930
transform 1 0 456 0 -1 770
box -8 -3 46 105
use NAND2X1  NAND2X1_67
timestamp 1681708930
transform -1 0 520 0 -1 770
box -8 -3 32 105
use XOR2X1  XOR2X1_150
timestamp 1681708930
transform -1 0 576 0 -1 770
box -8 -3 64 105
use FILL  FILL_1165
timestamp 1681708930
transform 1 0 576 0 -1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_106
timestamp 1681708930
transform -1 0 616 0 -1 770
box -8 -3 40 105
use FILL  FILL_1166
timestamp 1681708930
transform 1 0 616 0 -1 770
box -8 -3 16 105
use FILL  FILL_1171
timestamp 1681708930
transform 1 0 624 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_190
timestamp 1681708930
transform -1 0 648 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_191
timestamp 1681708930
transform -1 0 664 0 -1 770
box -9 -3 26 105
use FILL  FILL_1172
timestamp 1681708930
transform 1 0 664 0 -1 770
box -8 -3 16 105
use FILL  FILL_1174
timestamp 1681708930
transform 1 0 672 0 -1 770
box -8 -3 16 105
use FILL  FILL_1175
timestamp 1681708930
transform 1 0 680 0 -1 770
box -8 -3 16 105
use XOR2X1  XOR2X1_151
timestamp 1681708930
transform 1 0 688 0 -1 770
box -8 -3 64 105
use FILL  FILL_1176
timestamp 1681708930
transform 1 0 744 0 -1 770
box -8 -3 16 105
use FILL  FILL_1179
timestamp 1681708930
transform 1 0 752 0 -1 770
box -8 -3 16 105
use FILL  FILL_1180
timestamp 1681708930
transform 1 0 760 0 -1 770
box -8 -3 16 105
use FILL  FILL_1181
timestamp 1681708930
transform 1 0 768 0 -1 770
box -8 -3 16 105
use FILL  FILL_1182
timestamp 1681708930
transform 1 0 776 0 -1 770
box -8 -3 16 105
use FILL  FILL_1183
timestamp 1681708930
transform 1 0 784 0 -1 770
box -8 -3 16 105
use FILL  FILL_1184
timestamp 1681708930
transform 1 0 792 0 -1 770
box -8 -3 16 105
use FILL  FILL_1185
timestamp 1681708930
transform 1 0 800 0 -1 770
box -8 -3 16 105
use FILL  FILL_1186
timestamp 1681708930
transform 1 0 808 0 -1 770
box -8 -3 16 105
use FILL  FILL_1187
timestamp 1681708930
transform 1 0 816 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_68
timestamp 1681708930
transform -1 0 848 0 -1 770
box -8 -3 32 105
use FILL  FILL_1188
timestamp 1681708930
transform 1 0 848 0 -1 770
box -8 -3 16 105
use FILL  FILL_1190
timestamp 1681708930
transform 1 0 856 0 -1 770
box -8 -3 16 105
use FILL  FILL_1197
timestamp 1681708930
transform 1 0 864 0 -1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_110
timestamp 1681708930
transform 1 0 872 0 -1 770
box -8 -3 40 105
use FILL  FILL_1198
timestamp 1681708930
transform 1 0 904 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_193
timestamp 1681708930
transform -1 0 928 0 -1 770
box -9 -3 26 105
use FILL  FILL_1199
timestamp 1681708930
transform 1 0 928 0 -1 770
box -8 -3 16 105
use FILL  FILL_1200
timestamp 1681708930
transform 1 0 936 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_67
timestamp 1681708930
transform 1 0 944 0 -1 770
box -8 -3 46 105
use FILL  FILL_1201
timestamp 1681708930
transform 1 0 984 0 -1 770
box -8 -3 16 105
use FILL  FILL_1204
timestamp 1681708930
transform 1 0 992 0 -1 770
box -8 -3 16 105
use FILL  FILL_1205
timestamp 1681708930
transform 1 0 1000 0 -1 770
box -8 -3 16 105
use FILL  FILL_1206
timestamp 1681708930
transform 1 0 1008 0 -1 770
box -8 -3 16 105
use FILL  FILL_1207
timestamp 1681708930
transform 1 0 1016 0 -1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_111
timestamp 1681708930
transform -1 0 1056 0 -1 770
box -8 -3 40 105
use FILL  FILL_1208
timestamp 1681708930
transform 1 0 1056 0 -1 770
box -8 -3 16 105
use FILL  FILL_1209
timestamp 1681708930
transform 1 0 1064 0 -1 770
box -8 -3 16 105
use FILL  FILL_1210
timestamp 1681708930
transform 1 0 1072 0 -1 770
box -8 -3 16 105
use FILL  FILL_1217
timestamp 1681708930
transform 1 0 1080 0 -1 770
box -8 -3 16 105
use FILL  FILL_1218
timestamp 1681708930
transform 1 0 1088 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_196
timestamp 1681708930
transform -1 0 1112 0 -1 770
box -9 -3 26 105
use FILL  FILL_1219
timestamp 1681708930
transform 1 0 1112 0 -1 770
box -8 -3 16 105
use FILL  FILL_1220
timestamp 1681708930
transform 1 0 1120 0 -1 770
box -8 -3 16 105
use FILL  FILL_1221
timestamp 1681708930
transform 1 0 1128 0 -1 770
box -8 -3 16 105
use FILL  FILL_1222
timestamp 1681708930
transform 1 0 1136 0 -1 770
box -8 -3 16 105
use XOR2X1  XOR2X1_158
timestamp 1681708930
transform -1 0 1200 0 -1 770
box -8 -3 64 105
use XOR2X1  XOR2X1_159
timestamp 1681708930
transform -1 0 1256 0 -1 770
box -8 -3 64 105
use XOR2X1  XOR2X1_160
timestamp 1681708930
transform 1 0 1256 0 -1 770
box -8 -3 64 105
use XOR2X1  XOR2X1_161
timestamp 1681708930
transform -1 0 1368 0 -1 770
box -8 -3 64 105
use XOR2X1  XOR2X1_162
timestamp 1681708930
transform 1 0 1368 0 -1 770
box -8 -3 64 105
use XOR2X1  XOR2X1_163
timestamp 1681708930
transform -1 0 1480 0 -1 770
box -8 -3 64 105
use FILL  FILL_1223
timestamp 1681708930
transform 1 0 1480 0 -1 770
box -8 -3 16 105
use FILL  FILL_1224
timestamp 1681708930
transform 1 0 1488 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_26
timestamp 1681708930
transform 1 0 1496 0 -1 770
box -8 -3 46 105
use INVX2  INVX2_197
timestamp 1681708930
transform 1 0 1536 0 -1 770
box -9 -3 26 105
use FILL  FILL_1225
timestamp 1681708930
transform 1 0 1552 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_70
timestamp 1681708930
transform 1 0 1560 0 -1 770
box -8 -3 46 105
use FILL  FILL_1226
timestamp 1681708930
transform 1 0 1600 0 -1 770
box -8 -3 16 105
use FILL  FILL_1227
timestamp 1681708930
transform 1 0 1608 0 -1 770
box -8 -3 16 105
use FILL  FILL_1228
timestamp 1681708930
transform 1 0 1616 0 -1 770
box -8 -3 16 105
use FILL  FILL_1229
timestamp 1681708930
transform 1 0 1624 0 -1 770
box -8 -3 16 105
use FILL  FILL_1230
timestamp 1681708930
transform 1 0 1632 0 -1 770
box -8 -3 16 105
use FILL  FILL_1231
timestamp 1681708930
transform 1 0 1640 0 -1 770
box -8 -3 16 105
use FILL  FILL_1232
timestamp 1681708930
transform 1 0 1648 0 -1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_114
timestamp 1681708930
transform 1 0 1656 0 -1 770
box -8 -3 40 105
use FILL  FILL_1246
timestamp 1681708930
transform 1 0 1688 0 -1 770
box -8 -3 16 105
use FILL  FILL_1247
timestamp 1681708930
transform 1 0 1696 0 -1 770
box -8 -3 16 105
use FILL  FILL_1248
timestamp 1681708930
transform 1 0 1704 0 -1 770
box -8 -3 16 105
use BUFX2  BUFX2_8
timestamp 1681708930
transform 1 0 1712 0 -1 770
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_72
timestamp 1681708930
transform -1 0 1832 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_201
timestamp 1681708930
transform -1 0 1848 0 -1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_73
timestamp 1681708930
transform -1 0 1944 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_202
timestamp 1681708930
transform 1 0 1944 0 -1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_74
timestamp 1681708930
transform -1 0 2056 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_75
timestamp 1681708930
transform -1 0 2152 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_203
timestamp 1681708930
transform -1 0 2168 0 -1 770
box -9 -3 26 105
use FILL  FILL_1249
timestamp 1681708930
transform 1 0 2168 0 -1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_115
timestamp 1681708930
transform 1 0 2176 0 -1 770
box -8 -3 40 105
use FILL  FILL_1252
timestamp 1681708930
transform 1 0 2208 0 -1 770
box -8 -3 16 105
use FILL  FILL_1253
timestamp 1681708930
transform 1 0 2216 0 -1 770
box -8 -3 16 105
use FILL  FILL_1254
timestamp 1681708930
transform 1 0 2224 0 -1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_117
timestamp 1681708930
transform 1 0 2232 0 -1 770
box -8 -3 40 105
use NOR2X1  NOR2X1_66
timestamp 1681708930
transform -1 0 2288 0 -1 770
box -8 -3 32 105
use FILL  FILL_1269
timestamp 1681708930
transform 1 0 2288 0 -1 770
box -8 -3 16 105
use FILL  FILL_1270
timestamp 1681708930
transform 1 0 2296 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_207
timestamp 1681708930
transform 1 0 2304 0 -1 770
box -9 -3 26 105
use NAND2X1  NAND2X1_73
timestamp 1681708930
transform 1 0 2320 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_74
timestamp 1681708930
transform 1 0 2344 0 -1 770
box -8 -3 32 105
use FILL  FILL_1271
timestamp 1681708930
transform 1 0 2368 0 -1 770
box -8 -3 16 105
use FILL  FILL_1272
timestamp 1681708930
transform 1 0 2376 0 -1 770
box -8 -3 16 105
use FILL  FILL_1273
timestamp 1681708930
transform 1 0 2384 0 -1 770
box -8 -3 16 105
use FILL  FILL_1274
timestamp 1681708930
transform 1 0 2392 0 -1 770
box -8 -3 16 105
use FILL  FILL_1275
timestamp 1681708930
transform 1 0 2400 0 -1 770
box -8 -3 16 105
use FILL  FILL_1276
timestamp 1681708930
transform 1 0 2408 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_75
timestamp 1681708930
transform 1 0 2416 0 -1 770
box -8 -3 32 105
use XOR2X1  XOR2X1_167
timestamp 1681708930
transform -1 0 2496 0 -1 770
box -8 -3 64 105
use NAND3X1  NAND3X1_118
timestamp 1681708930
transform 1 0 2496 0 -1 770
box -8 -3 40 105
use XOR2X1  XOR2X1_168
timestamp 1681708930
transform -1 0 2584 0 -1 770
box -8 -3 64 105
use INVX2  INVX2_208
timestamp 1681708930
transform 1 0 2584 0 -1 770
box -9 -3 26 105
use XOR2X1  XOR2X1_169
timestamp 1681708930
transform -1 0 2656 0 -1 770
box -8 -3 64 105
use FILL  FILL_1277
timestamp 1681708930
transform 1 0 2656 0 -1 770
box -8 -3 16 105
use top_mod_new_VIA0  top_mod_new_VIA0_39
timestamp 1681708930
transform 1 0 2712 0 1 670
box -10 -3 10 3
use M3_M2  M3_M2_3072
timestamp 1681708930
transform 1 0 76 0 1 665
box -3 -3 3 3
use M2_M1  M2_M1_3154
timestamp 1681708930
transform 1 0 76 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3135
timestamp 1681708930
transform 1 0 84 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_3155
timestamp 1681708930
transform 1 0 132 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3157
timestamp 1681708930
transform 1 0 132 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_3223
timestamp 1681708930
transform 1 0 156 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3207
timestamp 1681708930
transform 1 0 156 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3077
timestamp 1681708930
transform 1 0 180 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3078
timestamp 1681708930
transform 1 0 236 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3136
timestamp 1681708930
transform 1 0 220 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3096
timestamp 1681708930
transform 1 0 292 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3108
timestamp 1681708930
transform 1 0 276 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_3137
timestamp 1681708930
transform 1 0 292 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3156
timestamp 1681708930
transform 1 0 228 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3157
timestamp 1681708930
transform 1 0 260 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3158
timestamp 1681708930
transform 1 0 276 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3224
timestamp 1681708930
transform 1 0 180 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3158
timestamp 1681708930
transform 1 0 204 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_3225
timestamp 1681708930
transform 1 0 268 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3175
timestamp 1681708930
transform 1 0 228 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3109
timestamp 1681708930
transform 1 0 332 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_3138
timestamp 1681708930
transform 1 0 396 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3159
timestamp 1681708930
transform 1 0 300 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3160
timestamp 1681708930
transform 1 0 356 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3226
timestamp 1681708930
transform 1 0 292 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3227
timestamp 1681708930
transform 1 0 380 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3228
timestamp 1681708930
transform 1 0 396 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3137
timestamp 1681708930
transform 1 0 420 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3138
timestamp 1681708930
transform 1 0 444 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3079
timestamp 1681708930
transform 1 0 492 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3085
timestamp 1681708930
transform 1 0 508 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3097
timestamp 1681708930
transform 1 0 492 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_3139
timestamp 1681708930
transform 1 0 468 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3161
timestamp 1681708930
transform 1 0 452 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3229
timestamp 1681708930
transform 1 0 420 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3230
timestamp 1681708930
transform 1 0 428 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3176
timestamp 1681708930
transform 1 0 292 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3177
timestamp 1681708930
transform 1 0 356 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3178
timestamp 1681708930
transform 1 0 396 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3179
timestamp 1681708930
transform 1 0 412 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3208
timestamp 1681708930
transform 1 0 380 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3209
timestamp 1681708930
transform 1 0 444 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_3140
timestamp 1681708930
transform 1 0 612 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3162
timestamp 1681708930
transform 1 0 476 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3163
timestamp 1681708930
transform 1 0 492 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3164
timestamp 1681708930
transform 1 0 508 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3165
timestamp 1681708930
transform 1 0 516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3166
timestamp 1681708930
transform 1 0 572 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3231
timestamp 1681708930
transform 1 0 468 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3232
timestamp 1681708930
transform 1 0 484 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3233
timestamp 1681708930
transform 1 0 500 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3180
timestamp 1681708930
transform 1 0 500 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3139
timestamp 1681708930
transform 1 0 596 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_3234
timestamp 1681708930
transform 1 0 596 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3235
timestamp 1681708930
transform 1 0 612 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3181
timestamp 1681708930
transform 1 0 572 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3182
timestamp 1681708930
transform 1 0 612 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3210
timestamp 1681708930
transform 1 0 484 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3211
timestamp 1681708930
transform 1 0 508 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3212
timestamp 1681708930
transform 1 0 580 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3110
timestamp 1681708930
transform 1 0 636 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_3141
timestamp 1681708930
transform 1 0 668 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3167
timestamp 1681708930
transform 1 0 644 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3168
timestamp 1681708930
transform 1 0 652 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3236
timestamp 1681708930
transform 1 0 636 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3213
timestamp 1681708930
transform 1 0 628 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_3169
timestamp 1681708930
transform 1 0 676 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3170
timestamp 1681708930
transform 1 0 708 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3140
timestamp 1681708930
transform 1 0 756 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3080
timestamp 1681708930
transform 1 0 780 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_3171
timestamp 1681708930
transform 1 0 772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3237
timestamp 1681708930
transform 1 0 668 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3159
timestamp 1681708930
transform 1 0 676 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3160
timestamp 1681708930
transform 1 0 708 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_3238
timestamp 1681708930
transform 1 0 756 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3214
timestamp 1681708930
transform 1 0 660 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3183
timestamp 1681708930
transform 1 0 692 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3184
timestamp 1681708930
transform 1 0 740 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3098
timestamp 1681708930
transform 1 0 852 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3111
timestamp 1681708930
transform 1 0 820 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3099
timestamp 1681708930
transform 1 0 892 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3112
timestamp 1681708930
transform 1 0 876 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_3172
timestamp 1681708930
transform 1 0 820 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3173
timestamp 1681708930
transform 1 0 852 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3174
timestamp 1681708930
transform 1 0 876 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3175
timestamp 1681708930
transform 1 0 892 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3239
timestamp 1681708930
transform 1 0 788 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3240
timestamp 1681708930
transform 1 0 796 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3241
timestamp 1681708930
transform 1 0 844 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3242
timestamp 1681708930
transform 1 0 852 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3243
timestamp 1681708930
transform 1 0 868 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3161
timestamp 1681708930
transform 1 0 876 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_3244
timestamp 1681708930
transform 1 0 884 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3185
timestamp 1681708930
transform 1 0 844 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3186
timestamp 1681708930
transform 1 0 868 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3187
timestamp 1681708930
transform 1 0 884 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3215
timestamp 1681708930
transform 1 0 804 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3216
timestamp 1681708930
transform 1 0 836 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3217
timestamp 1681708930
transform 1 0 860 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3113
timestamp 1681708930
transform 1 0 908 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3141
timestamp 1681708930
transform 1 0 900 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_3245
timestamp 1681708930
transform 1 0 900 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3246
timestamp 1681708930
transform 1 0 908 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3300
timestamp 1681708930
transform 1 0 908 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3176
timestamp 1681708930
transform 1 0 924 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3177
timestamp 1681708930
transform 1 0 932 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3178
timestamp 1681708930
transform 1 0 948 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3247
timestamp 1681708930
transform 1 0 956 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3188
timestamp 1681708930
transform 1 0 932 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3114
timestamp 1681708930
transform 1 0 1004 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_3179
timestamp 1681708930
transform 1 0 980 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3180
timestamp 1681708930
transform 1 0 1020 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3115
timestamp 1681708930
transform 1 0 1036 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3116
timestamp 1681708930
transform 1 0 1068 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_3181
timestamp 1681708930
transform 1 0 1036 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3182
timestamp 1681708930
transform 1 0 1068 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3248
timestamp 1681708930
transform 1 0 988 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3249
timestamp 1681708930
transform 1 0 1004 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3250
timestamp 1681708930
transform 1 0 1012 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3251
timestamp 1681708930
transform 1 0 1028 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3252
timestamp 1681708930
transform 1 0 1044 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3189
timestamp 1681708930
transform 1 0 980 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_3301
timestamp 1681708930
transform 1 0 988 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3302
timestamp 1681708930
transform 1 0 1020 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_3117
timestamp 1681708930
transform 1 0 1116 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_3253
timestamp 1681708930
transform 1 0 1100 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3254
timestamp 1681708930
transform 1 0 1108 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3190
timestamp 1681708930
transform 1 0 1100 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3162
timestamp 1681708930
transform 1 0 1132 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3142
timestamp 1681708930
transform 1 0 1148 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_3183
timestamp 1681708930
transform 1 0 1156 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3184
timestamp 1681708930
transform 1 0 1172 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3255
timestamp 1681708930
transform 1 0 1148 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3163
timestamp 1681708930
transform 1 0 1164 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3086
timestamp 1681708930
transform 1 0 1196 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3118
timestamp 1681708930
transform 1 0 1188 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_3185
timestamp 1681708930
transform 1 0 1188 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3256
timestamp 1681708930
transform 1 0 1180 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3164
timestamp 1681708930
transform 1 0 1188 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3191
timestamp 1681708930
transform 1 0 1188 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_3186
timestamp 1681708930
transform 1 0 1212 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3303
timestamp 1681708930
transform 1 0 1212 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_3119
timestamp 1681708930
transform 1 0 1236 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3143
timestamp 1681708930
transform 1 0 1228 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_3257
timestamp 1681708930
transform 1 0 1228 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3258
timestamp 1681708930
transform 1 0 1236 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3192
timestamp 1681708930
transform 1 0 1228 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_3142
timestamp 1681708930
transform 1 0 1268 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3187
timestamp 1681708930
transform 1 0 1244 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3188
timestamp 1681708930
transform 1 0 1260 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3189
timestamp 1681708930
transform 1 0 1268 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3120
timestamp 1681708930
transform 1 0 1284 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3193
timestamp 1681708930
transform 1 0 1276 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3121
timestamp 1681708930
transform 1 0 1308 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_3259
timestamp 1681708930
transform 1 0 1300 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3122
timestamp 1681708930
transform 1 0 1364 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_3190
timestamp 1681708930
transform 1 0 1364 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3260
timestamp 1681708930
transform 1 0 1356 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3261
timestamp 1681708930
transform 1 0 1372 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3144
timestamp 1681708930
transform 1 0 1428 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3100
timestamp 1681708930
transform 1 0 1452 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_3262
timestamp 1681708930
transform 1 0 1420 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3263
timestamp 1681708930
transform 1 0 1428 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3264
timestamp 1681708930
transform 1 0 1444 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3143
timestamp 1681708930
transform 1 0 1452 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3191
timestamp 1681708930
transform 1 0 1452 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3194
timestamp 1681708930
transform 1 0 1420 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3195
timestamp 1681708930
transform 1 0 1444 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3081
timestamp 1681708930
transform 1 0 1476 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_3192
timestamp 1681708930
transform 1 0 1476 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3165
timestamp 1681708930
transform 1 0 1468 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_3265
timestamp 1681708930
transform 1 0 1476 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3087
timestamp 1681708930
transform 1 0 1500 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_3135
timestamp 1681708930
transform 1 0 1508 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_3144
timestamp 1681708930
transform 1 0 1492 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_3123
timestamp 1681708930
transform 1 0 1508 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_3145
timestamp 1681708930
transform 1 0 1516 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3193
timestamp 1681708930
transform 1 0 1500 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3166
timestamp 1681708930
transform 1 0 1492 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3167
timestamp 1681708930
transform 1 0 1524 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3073
timestamp 1681708930
transform 1 0 1540 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3124
timestamp 1681708930
transform 1 0 1548 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_3194
timestamp 1681708930
transform 1 0 1540 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3195
timestamp 1681708930
transform 1 0 1548 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3266
timestamp 1681708930
transform 1 0 1532 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3267
timestamp 1681708930
transform 1 0 1548 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3304
timestamp 1681708930
transform 1 0 1524 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_3074
timestamp 1681708930
transform 1 0 1564 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3082
timestamp 1681708930
transform 1 0 1564 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_3146
timestamp 1681708930
transform 1 0 1564 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_3145
timestamp 1681708930
transform 1 0 1564 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_3268
timestamp 1681708930
transform 1 0 1564 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3088
timestamp 1681708930
transform 1 0 1588 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_3147
timestamp 1681708930
transform 1 0 1588 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_3125
timestamp 1681708930
transform 1 0 1596 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_3196
timestamp 1681708930
transform 1 0 1588 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3089
timestamp 1681708930
transform 1 0 1652 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3101
timestamp 1681708930
transform 1 0 1628 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_3197
timestamp 1681708930
transform 1 0 1604 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3146
timestamp 1681708930
transform 1 0 1612 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_3198
timestamp 1681708930
transform 1 0 1628 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3147
timestamp 1681708930
transform 1 0 1636 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_3199
timestamp 1681708930
transform 1 0 1652 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3168
timestamp 1681708930
transform 1 0 1588 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_3269
timestamp 1681708930
transform 1 0 1596 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3169
timestamp 1681708930
transform 1 0 1604 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_3270
timestamp 1681708930
transform 1 0 1612 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3271
timestamp 1681708930
transform 1 0 1636 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3272
timestamp 1681708930
transform 1 0 1644 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3170
timestamp 1681708930
transform 1 0 1652 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3075
timestamp 1681708930
transform 1 0 1676 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3083
timestamp 1681708930
transform 1 0 1668 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_3200
timestamp 1681708930
transform 1 0 1660 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3273
timestamp 1681708930
transform 1 0 1660 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3171
timestamp 1681708930
transform 1 0 1668 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3084
timestamp 1681708930
transform 1 0 1692 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_3201
timestamp 1681708930
transform 1 0 1692 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3274
timestamp 1681708930
transform 1 0 1684 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3275
timestamp 1681708930
transform 1 0 1692 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3196
timestamp 1681708930
transform 1 0 1660 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_3305
timestamp 1681708930
transform 1 0 1668 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_3197
timestamp 1681708930
transform 1 0 1684 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_3306
timestamp 1681708930
transform 1 0 1700 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_3218
timestamp 1681708930
transform 1 0 1668 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3219
timestamp 1681708930
transform 1 0 1692 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3076
timestamp 1681708930
transform 1 0 1724 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3090
timestamp 1681708930
transform 1 0 1828 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3091
timestamp 1681708930
transform 1 0 1844 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3126
timestamp 1681708930
transform 1 0 1876 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3127
timestamp 1681708930
transform 1 0 1900 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3128
timestamp 1681708930
transform 1 0 1924 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_3202
timestamp 1681708930
transform 1 0 1724 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3148
timestamp 1681708930
transform 1 0 1748 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3149
timestamp 1681708930
transform 1 0 1772 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_3203
timestamp 1681708930
transform 1 0 1780 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3150
timestamp 1681708930
transform 1 0 1788 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_3204
timestamp 1681708930
transform 1 0 1836 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3276
timestamp 1681708930
transform 1 0 1716 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3277
timestamp 1681708930
transform 1 0 1724 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3198
timestamp 1681708930
transform 1 0 1716 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3220
timestamp 1681708930
transform 1 0 1724 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_3278
timestamp 1681708930
transform 1 0 1772 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3279
timestamp 1681708930
transform 1 0 1860 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3199
timestamp 1681708930
transform 1 0 1844 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_3205
timestamp 1681708930
transform 1 0 1892 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3206
timestamp 1681708930
transform 1 0 1900 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3207
timestamp 1681708930
transform 1 0 1932 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3280
timestamp 1681708930
transform 1 0 1924 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3129
timestamp 1681708930
transform 1 0 2020 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3151
timestamp 1681708930
transform 1 0 1964 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3152
timestamp 1681708930
transform 1 0 1988 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_3208
timestamp 1681708930
transform 1 0 2020 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3281
timestamp 1681708930
transform 1 0 1940 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3200
timestamp 1681708930
transform 1 0 1932 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_3282
timestamp 1681708930
transform 1 0 1996 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3201
timestamp 1681708930
transform 1 0 1996 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_3307
timestamp 1681708930
transform 1 0 2108 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_3102
timestamp 1681708930
transform 1 0 2124 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_3148
timestamp 1681708930
transform 1 0 2124 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3149
timestamp 1681708930
transform 1 0 2156 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3209
timestamp 1681708930
transform 1 0 2172 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3283
timestamp 1681708930
transform 1 0 2164 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3284
timestamp 1681708930
transform 1 0 2180 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3103
timestamp 1681708930
transform 1 0 2204 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_3150
timestamp 1681708930
transform 1 0 2196 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_3153
timestamp 1681708930
transform 1 0 2196 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3130
timestamp 1681708930
transform 1 0 2228 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3092
timestamp 1681708930
transform 1 0 2236 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3093
timestamp 1681708930
transform 1 0 2284 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3104
timestamp 1681708930
transform 1 0 2276 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_3210
timestamp 1681708930
transform 1 0 2236 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3211
timestamp 1681708930
transform 1 0 2244 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3154
timestamp 1681708930
transform 1 0 2252 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_3212
timestamp 1681708930
transform 1 0 2268 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3285
timestamp 1681708930
transform 1 0 2252 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3308
timestamp 1681708930
transform 1 0 2276 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3213
timestamp 1681708930
transform 1 0 2292 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3214
timestamp 1681708930
transform 1 0 2308 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3131
timestamp 1681708930
transform 1 0 2324 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_3286
timestamp 1681708930
transform 1 0 2324 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3215
timestamp 1681708930
transform 1 0 2356 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3151
timestamp 1681708930
transform 1 0 2420 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3287
timestamp 1681708930
transform 1 0 2412 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3221
timestamp 1681708930
transform 1 0 2396 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3172
timestamp 1681708930
transform 1 0 2420 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_3152
timestamp 1681708930
transform 1 0 2452 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3288
timestamp 1681708930
transform 1 0 2444 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3222
timestamp 1681708930
transform 1 0 2428 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3094
timestamp 1681708930
transform 1 0 2468 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_3136
timestamp 1681708930
transform 1 0 2468 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_3216
timestamp 1681708930
transform 1 0 2460 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3202
timestamp 1681708930
transform 1 0 2460 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3105
timestamp 1681708930
transform 1 0 2484 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3106
timestamp 1681708930
transform 1 0 2500 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3132
timestamp 1681708930
transform 1 0 2492 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_3153
timestamp 1681708930
transform 1 0 2500 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_3107
timestamp 1681708930
transform 1 0 2524 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3155
timestamp 1681708930
transform 1 0 2508 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3133
timestamp 1681708930
transform 1 0 2564 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3095
timestamp 1681708930
transform 1 0 2596 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_3217
timestamp 1681708930
transform 1 0 2524 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3218
timestamp 1681708930
transform 1 0 2548 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3219
timestamp 1681708930
transform 1 0 2564 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3289
timestamp 1681708930
transform 1 0 2492 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3290
timestamp 1681708930
transform 1 0 2500 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3223
timestamp 1681708930
transform 1 0 2484 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_3291
timestamp 1681708930
transform 1 0 2524 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3292
timestamp 1681708930
transform 1 0 2532 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3293
timestamp 1681708930
transform 1 0 2540 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3173
timestamp 1681708930
transform 1 0 2548 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3156
timestamp 1681708930
transform 1 0 2580 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_3220
timestamp 1681708930
transform 1 0 2596 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3294
timestamp 1681708930
transform 1 0 2564 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3295
timestamp 1681708930
transform 1 0 2572 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3296
timestamp 1681708930
transform 1 0 2580 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3297
timestamp 1681708930
transform 1 0 2596 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3203
timestamp 1681708930
transform 1 0 2532 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3204
timestamp 1681708930
transform 1 0 2548 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3205
timestamp 1681708930
transform 1 0 2564 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3224
timestamp 1681708930
transform 1 0 2524 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3174
timestamp 1681708930
transform 1 0 2604 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_3309
timestamp 1681708930
transform 1 0 2596 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3310
timestamp 1681708930
transform 1 0 2604 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_3225
timestamp 1681708930
transform 1 0 2580 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3134
timestamp 1681708930
transform 1 0 2636 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_3221
timestamp 1681708930
transform 1 0 2636 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3222
timestamp 1681708930
transform 1 0 2644 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3298
timestamp 1681708930
transform 1 0 2620 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3299
timestamp 1681708930
transform 1 0 2628 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3206
timestamp 1681708930
transform 1 0 2620 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3226
timestamp 1681708930
transform 1 0 2612 0 1 585
box -3 -3 3 3
use top_mod_new_VIA0  top_mod_new_VIA0_40
timestamp 1681708930
transform 1 0 48 0 1 570
box -10 -3 10 3
use M3_M2  M3_M2_3227
timestamp 1681708930
transform 1 0 84 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_76
timestamp 1681708930
transform -1 0 168 0 1 570
box -8 -3 104 105
use M3_M2  M3_M2_3228
timestamp 1681708930
transform 1 0 188 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_77
timestamp 1681708930
transform 1 0 168 0 1 570
box -8 -3 104 105
use OAI21X1  OAI21X1_75
timestamp 1681708930
transform 1 0 264 0 1 570
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_78
timestamp 1681708930
transform -1 0 392 0 1 570
box -8 -3 104 105
use OAI21X1  OAI21X1_76
timestamp 1681708930
transform -1 0 424 0 1 570
box -8 -3 34 105
use INVX2  INVX2_209
timestamp 1681708930
transform 1 0 424 0 1 570
box -9 -3 26 105
use M3_M2  M3_M2_3229
timestamp 1681708930
transform 1 0 460 0 1 575
box -3 -3 3 3
use OAI21X1  OAI21X1_77
timestamp 1681708930
transform 1 0 440 0 1 570
box -8 -3 34 105
use AOI22X1  AOI22X1_76
timestamp 1681708930
transform 1 0 472 0 1 570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_79
timestamp 1681708930
transform -1 0 608 0 1 570
box -8 -3 104 105
use OAI21X1  OAI21X1_78
timestamp 1681708930
transform -1 0 640 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_79
timestamp 1681708930
transform 1 0 640 0 1 570
box -8 -3 34 105
use M3_M2  M3_M2_3230
timestamp 1681708930
transform 1 0 772 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_80
timestamp 1681708930
transform -1 0 768 0 1 570
box -8 -3 104 105
use M3_M2  M3_M2_3231
timestamp 1681708930
transform 1 0 796 0 1 575
box -3 -3 3 3
use BUFX2  BUFX2_9
timestamp 1681708930
transform 1 0 768 0 1 570
box -5 -3 28 105
use M3_M2  M3_M2_3232
timestamp 1681708930
transform 1 0 852 0 1 575
box -3 -3 3 3
use XOR2X1  XOR2X1_170
timestamp 1681708930
transform -1 0 848 0 1 570
box -8 -3 64 105
use OAI22X1  OAI22X1_27
timestamp 1681708930
transform 1 0 848 0 1 570
box -8 -3 46 105
use INVX2  INVX2_210
timestamp 1681708930
transform -1 0 904 0 1 570
box -9 -3 26 105
use NOR2X1  NOR2X1_67
timestamp 1681708930
transform 1 0 904 0 1 570
box -8 -3 32 105
use AOI22X1  AOI22X1_77
timestamp 1681708930
transform 1 0 928 0 1 570
box -8 -3 46 105
use INVX2  INVX2_211
timestamp 1681708930
transform -1 0 984 0 1 570
box -9 -3 26 105
use M3_M2  M3_M2_3233
timestamp 1681708930
transform 1 0 1020 0 1 575
box -3 -3 3 3
use AOI21X1  AOI21X1_41
timestamp 1681708930
transform -1 0 1016 0 1 570
box -7 -3 39 105
use NOR2X1  NOR2X1_68
timestamp 1681708930
transform 1 0 1016 0 1 570
box -8 -3 32 105
use XOR2X1  XOR2X1_171
timestamp 1681708930
transform -1 0 1096 0 1 570
box -8 -3 64 105
use FILL  FILL_1278
timestamp 1681708930
transform 1 0 1096 0 1 570
box -8 -3 16 105
use INVX2  INVX2_212
timestamp 1681708930
transform 1 0 1104 0 1 570
box -9 -3 26 105
use FILL  FILL_1279
timestamp 1681708930
transform 1 0 1120 0 1 570
box -8 -3 16 105
use FILL  FILL_1280
timestamp 1681708930
transform 1 0 1128 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_78
timestamp 1681708930
transform -1 0 1176 0 1 570
box -8 -3 46 105
use FILL  FILL_1281
timestamp 1681708930
transform 1 0 1176 0 1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_69
timestamp 1681708930
transform -1 0 1208 0 1 570
box -8 -3 32 105
use FILL  FILL_1282
timestamp 1681708930
transform 1 0 1208 0 1 570
box -8 -3 16 105
use INVX2  INVX2_213
timestamp 1681708930
transform -1 0 1232 0 1 570
box -9 -3 26 105
use INVX2  INVX2_214
timestamp 1681708930
transform 1 0 1232 0 1 570
box -9 -3 26 105
use NAND2X1  NAND2X1_76
timestamp 1681708930
transform 1 0 1248 0 1 570
box -8 -3 32 105
use FILL  FILL_1283
timestamp 1681708930
transform 1 0 1272 0 1 570
box -8 -3 16 105
use FILL  FILL_1284
timestamp 1681708930
transform 1 0 1280 0 1 570
box -8 -3 16 105
use FILL  FILL_1285
timestamp 1681708930
transform 1 0 1288 0 1 570
box -8 -3 16 105
use FILL  FILL_1286
timestamp 1681708930
transform 1 0 1296 0 1 570
box -8 -3 16 105
use XNOR2X1  XNOR2X1_49
timestamp 1681708930
transform -1 0 1360 0 1 570
box -8 -3 64 105
use FILL  FILL_1287
timestamp 1681708930
transform 1 0 1360 0 1 570
box -8 -3 16 105
use XOR2X1  XOR2X1_172
timestamp 1681708930
transform -1 0 1424 0 1 570
box -8 -3 64 105
use INVX2  INVX2_215
timestamp 1681708930
transform 1 0 1424 0 1 570
box -9 -3 26 105
use FILL  FILL_1288
timestamp 1681708930
transform 1 0 1440 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_80
timestamp 1681708930
transform -1 0 1480 0 1 570
box -8 -3 34 105
use FILL  FILL_1289
timestamp 1681708930
transform 1 0 1480 0 1 570
box -8 -3 16 105
use NAND3X1  NAND3X1_119
timestamp 1681708930
transform 1 0 1488 0 1 570
box -8 -3 40 105
use NOR2X1  NOR2X1_70
timestamp 1681708930
transform 1 0 1520 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_77
timestamp 1681708930
transform 1 0 1544 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_78
timestamp 1681708930
transform 1 0 1568 0 1 570
box -8 -3 32 105
use INVX2  INVX2_216
timestamp 1681708930
transform 1 0 1592 0 1 570
box -9 -3 26 105
use AOI22X1  AOI22X1_79
timestamp 1681708930
transform -1 0 1648 0 1 570
box -8 -3 46 105
use INVX2  INVX2_217
timestamp 1681708930
transform -1 0 1664 0 1 570
box -9 -3 26 105
use AOI21X1  AOI21X1_42
timestamp 1681708930
transform -1 0 1696 0 1 570
box -7 -3 39 105
use NOR2X1  NOR2X1_71
timestamp 1681708930
transform 1 0 1696 0 1 570
box -8 -3 32 105
use M3_M2  M3_M2_3234
timestamp 1681708930
transform 1 0 1764 0 1 575
box -3 -3 3 3
use XOR2X1  XOR2X1_173
timestamp 1681708930
transform -1 0 1776 0 1 570
box -8 -3 64 105
use M3_M2  M3_M2_3235
timestamp 1681708930
transform 1 0 1788 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3236
timestamp 1681708930
transform 1 0 1828 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3237
timestamp 1681708930
transform 1 0 1852 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_81
timestamp 1681708930
transform -1 0 1872 0 1 570
box -8 -3 104 105
use XOR2X1  XOR2X1_174
timestamp 1681708930
transform -1 0 1928 0 1 570
box -8 -3 64 105
use FILL  FILL_1290
timestamp 1681708930
transform 1 0 1928 0 1 570
box -8 -3 16 105
use XOR2X1  XOR2X1_175
timestamp 1681708930
transform -1 0 1992 0 1 570
box -8 -3 64 105
use XOR2X1  XOR2X1_176
timestamp 1681708930
transform 1 0 1992 0 1 570
box -8 -3 64 105
use FILL  FILL_1291
timestamp 1681708930
transform 1 0 2048 0 1 570
box -8 -3 16 105
use FILL  FILL_1292
timestamp 1681708930
transform 1 0 2056 0 1 570
box -8 -3 16 105
use FILL  FILL_1293
timestamp 1681708930
transform 1 0 2064 0 1 570
box -8 -3 16 105
use OR2X1  OR2X1_21
timestamp 1681708930
transform -1 0 2104 0 1 570
box -8 -3 40 105
use FILL  FILL_1294
timestamp 1681708930
transform 1 0 2104 0 1 570
box -8 -3 16 105
use FILL  FILL_1295
timestamp 1681708930
transform 1 0 2112 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_81
timestamp 1681708930
transform -1 0 2152 0 1 570
box -8 -3 34 105
use FILL  FILL_1296
timestamp 1681708930
transform 1 0 2152 0 1 570
box -8 -3 16 105
use FILL  FILL_1323
timestamp 1681708930
transform 1 0 2160 0 1 570
box -8 -3 16 105
use FILL  FILL_1325
timestamp 1681708930
transform 1 0 2168 0 1 570
box -8 -3 16 105
use FILL  FILL_1327
timestamp 1681708930
transform 1 0 2176 0 1 570
box -8 -3 16 105
use FILL  FILL_1329
timestamp 1681708930
transform 1 0 2184 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_86
timestamp 1681708930
transform -1 0 2224 0 1 570
box -8 -3 34 105
use FILL  FILL_1330
timestamp 1681708930
transform 1 0 2224 0 1 570
box -8 -3 16 105
use FILL  FILL_1331
timestamp 1681708930
transform 1 0 2232 0 1 570
box -8 -3 16 105
use AOI21X1  AOI21X1_45
timestamp 1681708930
transform 1 0 2240 0 1 570
box -7 -3 39 105
use NOR2X1  NOR2X1_76
timestamp 1681708930
transform 1 0 2272 0 1 570
box -8 -3 32 105
use FILL  FILL_1332
timestamp 1681708930
transform 1 0 2296 0 1 570
box -8 -3 16 105
use INVX2  INVX2_228
timestamp 1681708930
transform 1 0 2304 0 1 570
box -9 -3 26 105
use FILL  FILL_1344
timestamp 1681708930
transform 1 0 2320 0 1 570
box -8 -3 16 105
use FILL  FILL_1348
timestamp 1681708930
transform 1 0 2328 0 1 570
box -8 -3 16 105
use FILL  FILL_1350
timestamp 1681708930
transform 1 0 2336 0 1 570
box -8 -3 16 105
use FILL  FILL_1352
timestamp 1681708930
transform 1 0 2344 0 1 570
box -8 -3 16 105
use FILL  FILL_1353
timestamp 1681708930
transform 1 0 2352 0 1 570
box -8 -3 16 105
use XNOR2X1  XNOR2X1_50
timestamp 1681708930
transform -1 0 2416 0 1 570
box -8 -3 64 105
use FILL  FILL_1354
timestamp 1681708930
transform 1 0 2416 0 1 570
box -8 -3 16 105
use NAND3X1  NAND3X1_126
timestamp 1681708930
transform -1 0 2456 0 1 570
box -8 -3 40 105
use FILL  FILL_1355
timestamp 1681708930
transform 1 0 2456 0 1 570
box -8 -3 16 105
use FILL  FILL_1356
timestamp 1681708930
transform 1 0 2464 0 1 570
box -8 -3 16 105
use FILL  FILL_1357
timestamp 1681708930
transform 1 0 2472 0 1 570
box -8 -3 16 105
use INVX2  INVX2_229
timestamp 1681708930
transform -1 0 2496 0 1 570
box -9 -3 26 105
use OAI21X1  OAI21X1_87
timestamp 1681708930
transform -1 0 2528 0 1 570
box -8 -3 34 105
use AOI22X1  AOI22X1_86
timestamp 1681708930
transform 1 0 2528 0 1 570
box -8 -3 46 105
use AOI21X1  AOI21X1_46
timestamp 1681708930
transform 1 0 2568 0 1 570
box -7 -3 39 105
use NOR2X1  NOR2X1_77
timestamp 1681708930
transform 1 0 2600 0 1 570
box -8 -3 32 105
use FILL  FILL_1358
timestamp 1681708930
transform 1 0 2624 0 1 570
box -8 -3 16 105
use INVX2  INVX2_230
timestamp 1681708930
transform 1 0 2632 0 1 570
box -9 -3 26 105
use FILL  FILL_1359
timestamp 1681708930
transform 1 0 2648 0 1 570
box -8 -3 16 105
use FILL  FILL_1372
timestamp 1681708930
transform 1 0 2656 0 1 570
box -8 -3 16 105
use top_mod_new_VIA0  top_mod_new_VIA0_41
timestamp 1681708930
transform 1 0 2688 0 1 570
box -10 -3 10 3
use M3_M2  M3_M2_3296
timestamp 1681708930
transform 1 0 68 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_3267
timestamp 1681708930
transform 1 0 148 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_3322
timestamp 1681708930
transform 1 0 172 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3323
timestamp 1681708930
transform 1 0 188 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3324
timestamp 1681708930
transform 1 0 204 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3395
timestamp 1681708930
transform 1 0 92 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3396
timestamp 1681708930
transform 1 0 148 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3325
timestamp 1681708930
transform 1 0 92 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_3464
timestamp 1681708930
transform 1 0 204 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3325
timestamp 1681708930
transform 1 0 236 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3326
timestamp 1681708930
transform 1 0 244 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_3326
timestamp 1681708930
transform 1 0 244 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3268
timestamp 1681708930
transform 1 0 284 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_3327
timestamp 1681708930
transform 1 0 284 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3328
timestamp 1681708930
transform 1 0 300 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3397
timestamp 1681708930
transform 1 0 268 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3305
timestamp 1681708930
transform 1 0 284 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_3398
timestamp 1681708930
transform 1 0 340 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3465
timestamp 1681708930
transform 1 0 284 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_3327
timestamp 1681708930
transform 1 0 324 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3238
timestamp 1681708930
transform 1 0 404 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3239
timestamp 1681708930
transform 1 0 428 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3269
timestamp 1681708930
transform 1 0 484 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3297
timestamp 1681708930
transform 1 0 452 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_3329
timestamp 1681708930
transform 1 0 484 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_3240
timestamp 1681708930
transform 1 0 524 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_3330
timestamp 1681708930
transform 1 0 508 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3331
timestamp 1681708930
transform 1 0 524 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_3241
timestamp 1681708930
transform 1 0 588 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3270
timestamp 1681708930
transform 1 0 548 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3271
timestamp 1681708930
transform 1 0 596 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3272
timestamp 1681708930
transform 1 0 660 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_3332
timestamp 1681708930
transform 1 0 548 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3333
timestamp 1681708930
transform 1 0 636 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_3298
timestamp 1681708930
transform 1 0 644 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_3334
timestamp 1681708930
transform 1 0 660 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3335
timestamp 1681708930
transform 1 0 668 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3399
timestamp 1681708930
transform 1 0 396 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3400
timestamp 1681708930
transform 1 0 404 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3401
timestamp 1681708930
transform 1 0 460 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3402
timestamp 1681708930
transform 1 0 500 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3403
timestamp 1681708930
transform 1 0 516 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3404
timestamp 1681708930
transform 1 0 532 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3405
timestamp 1681708930
transform 1 0 596 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3406
timestamp 1681708930
transform 1 0 628 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3407
timestamp 1681708930
transform 1 0 644 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3328
timestamp 1681708930
transform 1 0 484 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3329
timestamp 1681708930
transform 1 0 524 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3330
timestamp 1681708930
transform 1 0 580 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3373
timestamp 1681708930
transform 1 0 532 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3386
timestamp 1681708930
transform 1 0 604 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_3387
timestamp 1681708930
transform 1 0 636 0 1 485
box -3 -3 3 3
use M2_M1  M2_M1_3466
timestamp 1681708930
transform 1 0 668 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_3355
timestamp 1681708930
transform 1 0 668 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3388
timestamp 1681708930
transform 1 0 676 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_3273
timestamp 1681708930
transform 1 0 692 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_3336
timestamp 1681708930
transform 1 0 692 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_3242
timestamp 1681708930
transform 1 0 724 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_3337
timestamp 1681708930
transform 1 0 724 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3408
timestamp 1681708930
transform 1 0 692 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3409
timestamp 1681708930
transform 1 0 700 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3484
timestamp 1681708930
transform 1 0 692 0 1 505
box -2 -2 2 2
use M3_M2  M3_M2_3306
timestamp 1681708930
transform 1 0 708 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_3410
timestamp 1681708930
transform 1 0 716 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3411
timestamp 1681708930
transform 1 0 732 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3412
timestamp 1681708930
transform 1 0 740 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3331
timestamp 1681708930
transform 1 0 724 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3389
timestamp 1681708930
transform 1 0 700 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_3243
timestamp 1681708930
transform 1 0 780 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3252
timestamp 1681708930
transform 1 0 764 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3253
timestamp 1681708930
transform 1 0 788 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3274
timestamp 1681708930
transform 1 0 764 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3275
timestamp 1681708930
transform 1 0 804 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3276
timestamp 1681708930
transform 1 0 828 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_3338
timestamp 1681708930
transform 1 0 748 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3339
timestamp 1681708930
transform 1 0 756 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3340
timestamp 1681708930
transform 1 0 764 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3341
timestamp 1681708930
transform 1 0 780 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_3299
timestamp 1681708930
transform 1 0 788 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_3244
timestamp 1681708930
transform 1 0 876 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_3342
timestamp 1681708930
transform 1 0 796 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3343
timestamp 1681708930
transform 1 0 804 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3344
timestamp 1681708930
transform 1 0 820 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3345
timestamp 1681708930
transform 1 0 828 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3346
timestamp 1681708930
transform 1 0 844 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3347
timestamp 1681708930
transform 1 0 860 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3413
timestamp 1681708930
transform 1 0 772 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3414
timestamp 1681708930
transform 1 0 788 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3332
timestamp 1681708930
transform 1 0 780 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3307
timestamp 1681708930
transform 1 0 804 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_3415
timestamp 1681708930
transform 1 0 812 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3416
timestamp 1681708930
transform 1 0 828 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3417
timestamp 1681708930
transform 1 0 836 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3418
timestamp 1681708930
transform 1 0 852 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3333
timestamp 1681708930
transform 1 0 820 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3254
timestamp 1681708930
transform 1 0 964 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_3348
timestamp 1681708930
transform 1 0 924 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3349
timestamp 1681708930
transform 1 0 932 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3419
timestamp 1681708930
transform 1 0 892 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3420
timestamp 1681708930
transform 1 0 900 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3308
timestamp 1681708930
transform 1 0 932 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_3350
timestamp 1681708930
transform 1 0 980 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3421
timestamp 1681708930
transform 1 0 956 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3334
timestamp 1681708930
transform 1 0 860 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3335
timestamp 1681708930
transform 1 0 876 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3356
timestamp 1681708930
transform 1 0 852 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3357
timestamp 1681708930
transform 1 0 868 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3358
timestamp 1681708930
transform 1 0 908 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3336
timestamp 1681708930
transform 1 0 948 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3374
timestamp 1681708930
transform 1 0 900 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3375
timestamp 1681708930
transform 1 0 932 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3390
timestamp 1681708930
transform 1 0 924 0 1 485
box -3 -3 3 3
use M2_M1  M2_M1_3351
timestamp 1681708930
transform 1 0 1036 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3352
timestamp 1681708930
transform 1 0 1044 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3422
timestamp 1681708930
transform 1 0 1004 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3423
timestamp 1681708930
transform 1 0 1012 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3309
timestamp 1681708930
transform 1 0 1036 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_3245
timestamp 1681708930
transform 1 0 1092 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3255
timestamp 1681708930
transform 1 0 1092 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3277
timestamp 1681708930
transform 1 0 1108 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_3353
timestamp 1681708930
transform 1 0 1092 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3424
timestamp 1681708930
transform 1 0 1068 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3359
timestamp 1681708930
transform 1 0 1028 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3376
timestamp 1681708930
transform 1 0 1004 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3310
timestamp 1681708930
transform 1 0 1100 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_3300
timestamp 1681708930
transform 1 0 1124 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_3425
timestamp 1681708930
transform 1 0 1116 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3467
timestamp 1681708930
transform 1 0 1100 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_3278
timestamp 1681708930
transform 1 0 1140 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3301
timestamp 1681708930
transform 1 0 1156 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_3246
timestamp 1681708930
transform 1 0 1204 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3279
timestamp 1681708930
transform 1 0 1212 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_3354
timestamp 1681708930
transform 1 0 1172 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3355
timestamp 1681708930
transform 1 0 1188 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3356
timestamp 1681708930
transform 1 0 1204 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_3311
timestamp 1681708930
transform 1 0 1148 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_3426
timestamp 1681708930
transform 1 0 1156 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3468
timestamp 1681708930
transform 1 0 1132 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3469
timestamp 1681708930
transform 1 0 1140 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3485
timestamp 1681708930
transform 1 0 1124 0 1 505
box -2 -2 2 2
use M3_M2  M3_M2_3360
timestamp 1681708930
transform 1 0 1132 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3337
timestamp 1681708930
transform 1 0 1156 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_3427
timestamp 1681708930
transform 1 0 1180 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3470
timestamp 1681708930
transform 1 0 1164 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3486
timestamp 1681708930
transform 1 0 1148 0 1 505
box -2 -2 2 2
use M3_M2  M3_M2_3377
timestamp 1681708930
transform 1 0 1172 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_3428
timestamp 1681708930
transform 1 0 1212 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3338
timestamp 1681708930
transform 1 0 1204 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3247
timestamp 1681708930
transform 1 0 1268 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3280
timestamp 1681708930
transform 1 0 1244 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_3357
timestamp 1681708930
transform 1 0 1252 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3358
timestamp 1681708930
transform 1 0 1268 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3429
timestamp 1681708930
transform 1 0 1228 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3430
timestamp 1681708930
transform 1 0 1260 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3431
timestamp 1681708930
transform 1 0 1268 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3471
timestamp 1681708930
transform 1 0 1212 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3472
timestamp 1681708930
transform 1 0 1220 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_3339
timestamp 1681708930
transform 1 0 1228 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_3473
timestamp 1681708930
transform 1 0 1244 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_3340
timestamp 1681708930
transform 1 0 1252 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_3487
timestamp 1681708930
transform 1 0 1236 0 1 505
box -2 -2 2 2
use M3_M2  M3_M2_3361
timestamp 1681708930
transform 1 0 1244 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3302
timestamp 1681708930
transform 1 0 1292 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_3432
timestamp 1681708930
transform 1 0 1292 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3341
timestamp 1681708930
transform 1 0 1292 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3281
timestamp 1681708930
transform 1 0 1300 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_3311
timestamp 1681708930
transform 1 0 1308 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_3248
timestamp 1681708930
transform 1 0 1340 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_3312
timestamp 1681708930
transform 1 0 1340 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3359
timestamp 1681708930
transform 1 0 1300 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3360
timestamp 1681708930
transform 1 0 1324 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3361
timestamp 1681708930
transform 1 0 1332 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3433
timestamp 1681708930
transform 1 0 1300 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3312
timestamp 1681708930
transform 1 0 1324 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_3434
timestamp 1681708930
transform 1 0 1340 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3378
timestamp 1681708930
transform 1 0 1300 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3391
timestamp 1681708930
transform 1 0 1308 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_3256
timestamp 1681708930
transform 1 0 1364 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3282
timestamp 1681708930
transform 1 0 1356 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3283
timestamp 1681708930
transform 1 0 1380 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_3313
timestamp 1681708930
transform 1 0 1388 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3362
timestamp 1681708930
transform 1 0 1356 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3363
timestamp 1681708930
transform 1 0 1380 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_3313
timestamp 1681708930
transform 1 0 1356 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_3435
timestamp 1681708930
transform 1 0 1364 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3436
timestamp 1681708930
transform 1 0 1396 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3257
timestamp 1681708930
transform 1 0 1412 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_3314
timestamp 1681708930
transform 1 0 1412 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_3284
timestamp 1681708930
transform 1 0 1436 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_3364
timestamp 1681708930
transform 1 0 1428 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3365
timestamp 1681708930
transform 1 0 1436 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3437
timestamp 1681708930
transform 1 0 1412 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3438
timestamp 1681708930
transform 1 0 1436 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3314
timestamp 1681708930
transform 1 0 1444 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_3474
timestamp 1681708930
transform 1 0 1444 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_3362
timestamp 1681708930
transform 1 0 1428 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3258
timestamp 1681708930
transform 1 0 1484 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_3315
timestamp 1681708930
transform 1 0 1476 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3366
timestamp 1681708930
transform 1 0 1468 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3367
timestamp 1681708930
transform 1 0 1484 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3439
timestamp 1681708930
transform 1 0 1468 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3315
timestamp 1681708930
transform 1 0 1476 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_3342
timestamp 1681708930
transform 1 0 1468 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3392
timestamp 1681708930
transform 1 0 1460 0 1 485
box -3 -3 3 3
use M2_M1  M2_M1_3440
timestamp 1681708930
transform 1 0 1492 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3316
timestamp 1681708930
transform 1 0 1500 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_3368
timestamp 1681708930
transform 1 0 1532 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3441
timestamp 1681708930
transform 1 0 1516 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3442
timestamp 1681708930
transform 1 0 1532 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3475
timestamp 1681708930
transform 1 0 1500 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3476
timestamp 1681708930
transform 1 0 1516 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3488
timestamp 1681708930
transform 1 0 1508 0 1 505
box -2 -2 2 2
use M3_M2  M3_M2_3379
timestamp 1681708930
transform 1 0 1492 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3363
timestamp 1681708930
transform 1 0 1532 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3393
timestamp 1681708930
transform 1 0 1516 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_3285
timestamp 1681708930
transform 1 0 1580 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_3369
timestamp 1681708930
transform 1 0 1556 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_3303
timestamp 1681708930
transform 1 0 1564 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_3370
timestamp 1681708930
transform 1 0 1580 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_3304
timestamp 1681708930
transform 1 0 1588 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_3371
timestamp 1681708930
transform 1 0 1596 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3443
timestamp 1681708930
transform 1 0 1564 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3444
timestamp 1681708930
transform 1 0 1580 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3445
timestamp 1681708930
transform 1 0 1588 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3343
timestamp 1681708930
transform 1 0 1564 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3344
timestamp 1681708930
transform 1 0 1580 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3364
timestamp 1681708930
transform 1 0 1572 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3365
timestamp 1681708930
transform 1 0 1596 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3394
timestamp 1681708930
transform 1 0 1596 0 1 485
box -3 -3 3 3
use M2_M1  M2_M1_3372
timestamp 1681708930
transform 1 0 1620 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3446
timestamp 1681708930
transform 1 0 1628 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3447
timestamp 1681708930
transform 1 0 1636 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3345
timestamp 1681708930
transform 1 0 1628 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3380
timestamp 1681708930
transform 1 0 1636 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3286
timestamp 1681708930
transform 1 0 1660 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_3316
timestamp 1681708930
transform 1 0 1668 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3373
timestamp 1681708930
transform 1 0 1660 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_3366
timestamp 1681708930
transform 1 0 1668 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3259
timestamp 1681708930
transform 1 0 1708 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3287
timestamp 1681708930
transform 1 0 1700 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_3374
timestamp 1681708930
transform 1 0 1692 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3375
timestamp 1681708930
transform 1 0 1700 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3448
timestamp 1681708930
transform 1 0 1684 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3346
timestamp 1681708930
transform 1 0 1684 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_3449
timestamp 1681708930
transform 1 0 1716 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3381
timestamp 1681708930
transform 1 0 1724 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3395
timestamp 1681708930
transform 1 0 1716 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_3249
timestamp 1681708930
transform 1 0 1788 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3288
timestamp 1681708930
transform 1 0 1780 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3347
timestamp 1681708930
transform 1 0 1772 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_3376
timestamp 1681708930
transform 1 0 1788 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3377
timestamp 1681708930
transform 1 0 1796 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_3250
timestamp 1681708930
transform 1 0 1940 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3260
timestamp 1681708930
transform 1 0 1876 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3261
timestamp 1681708930
transform 1 0 1900 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_3378
timestamp 1681708930
transform 1 0 1844 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3379
timestamp 1681708930
transform 1 0 1852 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3380
timestamp 1681708930
transform 1 0 1900 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3381
timestamp 1681708930
transform 1 0 1908 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3450
timestamp 1681708930
transform 1 0 1812 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3451
timestamp 1681708930
transform 1 0 1852 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3317
timestamp 1681708930
transform 1 0 1876 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_3452
timestamp 1681708930
transform 1 0 1900 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3348
timestamp 1681708930
transform 1 0 1900 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3367
timestamp 1681708930
transform 1 0 1900 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_3453
timestamp 1681708930
transform 1 0 1956 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3368
timestamp 1681708930
transform 1 0 1988 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3262
timestamp 1681708930
transform 1 0 2020 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3289
timestamp 1681708930
transform 1 0 2012 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_3382
timestamp 1681708930
transform 1 0 2012 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3383
timestamp 1681708930
transform 1 0 2020 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_3349
timestamp 1681708930
transform 1 0 2020 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3369
timestamp 1681708930
transform 1 0 2052 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3290
timestamp 1681708930
transform 1 0 2076 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3370
timestamp 1681708930
transform 1 0 2092 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3263
timestamp 1681708930
transform 1 0 2108 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3291
timestamp 1681708930
transform 1 0 2124 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_3384
timestamp 1681708930
transform 1 0 2100 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3385
timestamp 1681708930
transform 1 0 2108 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_3318
timestamp 1681708930
transform 1 0 2100 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_3350
timestamp 1681708930
transform 1 0 2100 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_3454
timestamp 1681708930
transform 1 0 2116 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3455
timestamp 1681708930
transform 1 0 2140 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3477
timestamp 1681708930
transform 1 0 2124 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_3351
timestamp 1681708930
transform 1 0 2140 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_3489
timestamp 1681708930
transform 1 0 2132 0 1 505
box -2 -2 2 2
use M3_M2  M3_M2_3319
timestamp 1681708930
transform 1 0 2188 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_3478
timestamp 1681708930
transform 1 0 2180 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3479
timestamp 1681708930
transform 1 0 2188 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_3251
timestamp 1681708930
transform 1 0 2260 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_3456
timestamp 1681708930
transform 1 0 2252 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3352
timestamp 1681708930
transform 1 0 2252 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3264
timestamp 1681708930
transform 1 0 2276 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_3317
timestamp 1681708930
transform 1 0 2276 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3480
timestamp 1681708930
transform 1 0 2268 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_3292
timestamp 1681708930
transform 1 0 2292 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3353
timestamp 1681708930
transform 1 0 2292 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_3490
timestamp 1681708930
transform 1 0 2300 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_3481
timestamp 1681708930
transform 1 0 2316 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3318
timestamp 1681708930
transform 1 0 2332 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_3265
timestamp 1681708930
transform 1 0 2356 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3266
timestamp 1681708930
transform 1 0 2380 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3293
timestamp 1681708930
transform 1 0 2372 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_3386
timestamp 1681708930
transform 1 0 2372 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3387
timestamp 1681708930
transform 1 0 2380 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_3320
timestamp 1681708930
transform 1 0 2372 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_3294
timestamp 1681708930
transform 1 0 2412 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_3319
timestamp 1681708930
transform 1 0 2420 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3388
timestamp 1681708930
transform 1 0 2404 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3457
timestamp 1681708930
transform 1 0 2420 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3389
timestamp 1681708930
transform 1 0 2444 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3390
timestamp 1681708930
transform 1 0 2460 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_3382
timestamp 1681708930
transform 1 0 2436 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3295
timestamp 1681708930
transform 1 0 2508 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_3391
timestamp 1681708930
transform 1 0 2508 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3458
timestamp 1681708930
transform 1 0 2468 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3459
timestamp 1681708930
transform 1 0 2492 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3482
timestamp 1681708930
transform 1 0 2476 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_3321
timestamp 1681708930
transform 1 0 2500 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_3460
timestamp 1681708930
transform 1 0 2508 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3483
timestamp 1681708930
transform 1 0 2500 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_3354
timestamp 1681708930
transform 1 0 2508 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_3491
timestamp 1681708930
transform 1 0 2492 0 1 505
box -2 -2 2 2
use M3_M2  M3_M2_3371
timestamp 1681708930
transform 1 0 2500 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3383
timestamp 1681708930
transform 1 0 2476 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3384
timestamp 1681708930
transform 1 0 2492 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_3320
timestamp 1681708930
transform 1 0 2524 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3461
timestamp 1681708930
transform 1 0 2524 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3372
timestamp 1681708930
transform 1 0 2524 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3385
timestamp 1681708930
transform 1 0 2516 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3322
timestamp 1681708930
transform 1 0 2540 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_3321
timestamp 1681708930
transform 1 0 2580 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3392
timestamp 1681708930
transform 1 0 2564 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3393
timestamp 1681708930
transform 1 0 2572 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3462
timestamp 1681708930
transform 1 0 2556 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3323
timestamp 1681708930
transform 1 0 2572 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_3394
timestamp 1681708930
transform 1 0 2644 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3463
timestamp 1681708930
transform 1 0 2612 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_3324
timestamp 1681708930
transform 1 0 2644 0 1 525
box -3 -3 3 3
use top_mod_new_VIA0  top_mod_new_VIA0_42
timestamp 1681708930
transform 1 0 24 0 1 470
box -10 -3 10 3
use FILL  FILL_1297
timestamp 1681708930
transform 1 0 72 0 -1 570
box -8 -3 16 105
use FILL  FILL_1298
timestamp 1681708930
transform 1 0 80 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_82
timestamp 1681708930
transform -1 0 184 0 -1 570
box -8 -3 104 105
use NAND2X1  NAND2X1_79
timestamp 1681708930
transform 1 0 184 0 -1 570
box -8 -3 32 105
use OAI21X1  OAI21X1_82
timestamp 1681708930
transform -1 0 240 0 -1 570
box -8 -3 34 105
use INVX2  INVX2_218
timestamp 1681708930
transform 1 0 240 0 -1 570
box -9 -3 26 105
use OAI21X1  OAI21X1_83
timestamp 1681708930
transform 1 0 256 0 -1 570
box -8 -3 34 105
use M3_M2  M3_M2_3396
timestamp 1681708930
transform 1 0 380 0 1 475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_83
timestamp 1681708930
transform 1 0 288 0 -1 570
box -8 -3 104 105
use INVX2  INVX2_219
timestamp 1681708930
transform 1 0 384 0 -1 570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_84
timestamp 1681708930
transform -1 0 496 0 -1 570
box -8 -3 104 105
use M3_M2  M3_M2_3397
timestamp 1681708930
transform 1 0 516 0 1 475
box -3 -3 3 3
use AOI22X1  AOI22X1_80
timestamp 1681708930
transform 1 0 496 0 -1 570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_85
timestamp 1681708930
transform 1 0 536 0 -1 570
box -8 -3 104 105
use OAI21X1  OAI21X1_84
timestamp 1681708930
transform 1 0 632 0 -1 570
box -8 -3 34 105
use NAND2X1  NAND2X1_80
timestamp 1681708930
transform 1 0 664 0 -1 570
box -8 -3 32 105
use FILL  FILL_1299
timestamp 1681708930
transform 1 0 688 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_81
timestamp 1681708930
transform 1 0 696 0 -1 570
box -8 -3 46 105
use INVX2  INVX2_220
timestamp 1681708930
transform -1 0 752 0 -1 570
box -9 -3 26 105
use AOI22X1  AOI22X1_82
timestamp 1681708930
transform 1 0 752 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_83
timestamp 1681708930
transform 1 0 792 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_84
timestamp 1681708930
transform 1 0 832 0 -1 570
box -8 -3 46 105
use M3_M2  M3_M2_3398
timestamp 1681708930
transform 1 0 892 0 1 475
box -3 -3 3 3
use XOR2X1  XOR2X1_177
timestamp 1681708930
transform -1 0 928 0 -1 570
box -8 -3 64 105
use XOR2X1  XOR2X1_178
timestamp 1681708930
transform -1 0 984 0 -1 570
box -8 -3 64 105
use M3_M2  M3_M2_3399
timestamp 1681708930
transform 1 0 1068 0 1 475
box -3 -3 3 3
use XOR2X1  XOR2X1_179
timestamp 1681708930
transform -1 0 1040 0 -1 570
box -8 -3 64 105
use XOR2X1  XOR2X1_180
timestamp 1681708930
transform 1 0 1040 0 -1 570
box -8 -3 64 105
use NAND3X1  NAND3X1_120
timestamp 1681708930
transform -1 0 1128 0 -1 570
box -8 -3 40 105
use FILL  FILL_1300
timestamp 1681708930
transform 1 0 1128 0 -1 570
box -8 -3 16 105
use NAND3X1  NAND3X1_121
timestamp 1681708930
transform -1 0 1168 0 -1 570
box -8 -3 40 105
use OAI22X1  OAI22X1_28
timestamp 1681708930
transform -1 0 1208 0 -1 570
box -8 -3 46 105
use FILL  FILL_1301
timestamp 1681708930
transform 1 0 1208 0 -1 570
box -8 -3 16 105
use NAND3X1  NAND3X1_122
timestamp 1681708930
transform 1 0 1216 0 -1 570
box -8 -3 40 105
use INVX2  INVX2_221
timestamp 1681708930
transform 1 0 1248 0 -1 570
box -9 -3 26 105
use NAND2X1  NAND2X1_81
timestamp 1681708930
transform 1 0 1264 0 -1 570
box -8 -3 32 105
use INVX2  INVX2_222
timestamp 1681708930
transform -1 0 1304 0 -1 570
box -9 -3 26 105
use AOI21X1  AOI21X1_43
timestamp 1681708930
transform -1 0 1336 0 -1 570
box -7 -3 39 105
use NOR2X1  NOR2X1_72
timestamp 1681708930
transform 1 0 1336 0 -1 570
box -8 -3 32 105
use OR2X1  OR2X1_22
timestamp 1681708930
transform -1 0 1392 0 -1 570
box -8 -3 40 105
use INVX2  INVX2_223
timestamp 1681708930
transform -1 0 1408 0 -1 570
box -9 -3 26 105
use AOI21X1  AOI21X1_44
timestamp 1681708930
transform -1 0 1440 0 -1 570
box -7 -3 39 105
use OAI21X1  OAI21X1_85
timestamp 1681708930
transform -1 0 1472 0 -1 570
box -8 -3 34 105
use NOR2X1  NOR2X1_73
timestamp 1681708930
transform 1 0 1472 0 -1 570
box -8 -3 32 105
use NAND3X1  NAND3X1_123
timestamp 1681708930
transform -1 0 1528 0 -1 570
box -8 -3 40 105
use INVX2  INVX2_224
timestamp 1681708930
transform 1 0 1528 0 -1 570
box -9 -3 26 105
use AOI22X1  AOI22X1_85
timestamp 1681708930
transform 1 0 1544 0 -1 570
box -8 -3 46 105
use FILL  FILL_1302
timestamp 1681708930
transform 1 0 1584 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_225
timestamp 1681708930
transform 1 0 1592 0 -1 570
box -9 -3 26 105
use NOR2X1  NOR2X1_74
timestamp 1681708930
transform 1 0 1608 0 -1 570
box -8 -3 32 105
use FILL  FILL_1303
timestamp 1681708930
transform 1 0 1632 0 -1 570
box -8 -3 16 105
use FILL  FILL_1304
timestamp 1681708930
transform 1 0 1640 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_226
timestamp 1681708930
transform -1 0 1664 0 -1 570
box -9 -3 26 105
use NOR2X1  NOR2X1_75
timestamp 1681708930
transform 1 0 1664 0 -1 570
box -8 -3 32 105
use FILL  FILL_1305
timestamp 1681708930
transform 1 0 1688 0 -1 570
box -8 -3 16 105
use XOR2X1  XOR2X1_181
timestamp 1681708930
transform -1 0 1752 0 -1 570
box -8 -3 64 105
use FILL  FILL_1306
timestamp 1681708930
transform 1 0 1752 0 -1 570
box -8 -3 16 105
use FILL  FILL_1307
timestamp 1681708930
transform 1 0 1760 0 -1 570
box -8 -3 16 105
use FILL  FILL_1308
timestamp 1681708930
transform 1 0 1768 0 -1 570
box -8 -3 16 105
use FILL  FILL_1309
timestamp 1681708930
transform 1 0 1776 0 -1 570
box -8 -3 16 105
use FILL  FILL_1310
timestamp 1681708930
transform 1 0 1784 0 -1 570
box -8 -3 16 105
use XOR2X1  XOR2X1_182
timestamp 1681708930
transform -1 0 1848 0 -1 570
box -8 -3 64 105
use XOR2X1  XOR2X1_183
timestamp 1681708930
transform -1 0 1904 0 -1 570
box -8 -3 64 105
use XOR2X1  XOR2X1_184
timestamp 1681708930
transform -1 0 1960 0 -1 570
box -8 -3 64 105
use FILL  FILL_1311
timestamp 1681708930
transform 1 0 1960 0 -1 570
box -8 -3 16 105
use FILL  FILL_1312
timestamp 1681708930
transform 1 0 1968 0 -1 570
box -8 -3 16 105
use FILL  FILL_1313
timestamp 1681708930
transform 1 0 1976 0 -1 570
box -8 -3 16 105
use FILL  FILL_1314
timestamp 1681708930
transform 1 0 1984 0 -1 570
box -8 -3 16 105
use FILL  FILL_1315
timestamp 1681708930
transform 1 0 1992 0 -1 570
box -8 -3 16 105
use FILL  FILL_1316
timestamp 1681708930
transform 1 0 2000 0 -1 570
box -8 -3 16 105
use FILL  FILL_1317
timestamp 1681708930
transform 1 0 2008 0 -1 570
box -8 -3 16 105
use XOR2X1  XOR2X1_185
timestamp 1681708930
transform -1 0 2072 0 -1 570
box -8 -3 64 105
use FILL  FILL_1318
timestamp 1681708930
transform 1 0 2072 0 -1 570
box -8 -3 16 105
use FILL  FILL_1319
timestamp 1681708930
transform 1 0 2080 0 -1 570
box -8 -3 16 105
use FILL  FILL_1320
timestamp 1681708930
transform 1 0 2088 0 -1 570
box -8 -3 16 105
use FILL  FILL_1321
timestamp 1681708930
transform 1 0 2096 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_227
timestamp 1681708930
transform 1 0 2104 0 -1 570
box -9 -3 26 105
use NAND3X1  NAND3X1_124
timestamp 1681708930
transform -1 0 2152 0 -1 570
box -8 -3 40 105
use FILL  FILL_1322
timestamp 1681708930
transform 1 0 2152 0 -1 570
box -8 -3 16 105
use FILL  FILL_1324
timestamp 1681708930
transform 1 0 2160 0 -1 570
box -8 -3 16 105
use FILL  FILL_1326
timestamp 1681708930
transform 1 0 2168 0 -1 570
box -8 -3 16 105
use FILL  FILL_1328
timestamp 1681708930
transform 1 0 2176 0 -1 570
box -8 -3 16 105
use FILL  FILL_1333
timestamp 1681708930
transform 1 0 2184 0 -1 570
box -8 -3 16 105
use FILL  FILL_1334
timestamp 1681708930
transform 1 0 2192 0 -1 570
box -8 -3 16 105
use FILL  FILL_1335
timestamp 1681708930
transform 1 0 2200 0 -1 570
box -8 -3 16 105
use FILL  FILL_1336
timestamp 1681708930
transform 1 0 2208 0 -1 570
box -8 -3 16 105
use FILL  FILL_1337
timestamp 1681708930
transform 1 0 2216 0 -1 570
box -8 -3 16 105
use FILL  FILL_1338
timestamp 1681708930
transform 1 0 2224 0 -1 570
box -8 -3 16 105
use NAND3X1  NAND3X1_125
timestamp 1681708930
transform -1 0 2264 0 -1 570
box -8 -3 40 105
use FILL  FILL_1339
timestamp 1681708930
transform 1 0 2264 0 -1 570
box -8 -3 16 105
use FILL  FILL_1340
timestamp 1681708930
transform 1 0 2272 0 -1 570
box -8 -3 16 105
use FILL  FILL_1341
timestamp 1681708930
transform 1 0 2280 0 -1 570
box -8 -3 16 105
use FILL  FILL_1342
timestamp 1681708930
transform 1 0 2288 0 -1 570
box -8 -3 16 105
use FILL  FILL_1343
timestamp 1681708930
transform 1 0 2296 0 -1 570
box -8 -3 16 105
use FILL  FILL_1345
timestamp 1681708930
transform 1 0 2304 0 -1 570
box -8 -3 16 105
use FILL  FILL_1346
timestamp 1681708930
transform 1 0 2312 0 -1 570
box -8 -3 16 105
use FILL  FILL_1347
timestamp 1681708930
transform 1 0 2320 0 -1 570
box -8 -3 16 105
use FILL  FILL_1349
timestamp 1681708930
transform 1 0 2328 0 -1 570
box -8 -3 16 105
use FILL  FILL_1351
timestamp 1681708930
transform 1 0 2336 0 -1 570
box -8 -3 16 105
use FILL  FILL_1360
timestamp 1681708930
transform 1 0 2344 0 -1 570
box -8 -3 16 105
use AOI21X1  AOI21X1_47
timestamp 1681708930
transform -1 0 2384 0 -1 570
box -7 -3 39 105
use FILL  FILL_1361
timestamp 1681708930
transform 1 0 2384 0 -1 570
box -8 -3 16 105
use FILL  FILL_1362
timestamp 1681708930
transform 1 0 2392 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_231
timestamp 1681708930
transform 1 0 2400 0 -1 570
box -9 -3 26 105
use FILL  FILL_1363
timestamp 1681708930
transform 1 0 2416 0 -1 570
box -8 -3 16 105
use FILL  FILL_1364
timestamp 1681708930
transform 1 0 2424 0 -1 570
box -8 -3 16 105
use FILL  FILL_1365
timestamp 1681708930
transform 1 0 2432 0 -1 570
box -8 -3 16 105
use AOI21X1  AOI21X1_48
timestamp 1681708930
transform -1 0 2472 0 -1 570
box -7 -3 39 105
use NAND3X1  NAND3X1_127
timestamp 1681708930
transform -1 0 2504 0 -1 570
box -8 -3 40 105
use NOR2X1  NOR2X1_78
timestamp 1681708930
transform -1 0 2528 0 -1 570
box -8 -3 32 105
use FILL  FILL_1366
timestamp 1681708930
transform 1 0 2528 0 -1 570
box -8 -3 16 105
use FILL  FILL_1367
timestamp 1681708930
transform 1 0 2536 0 -1 570
box -8 -3 16 105
use FILL  FILL_1368
timestamp 1681708930
transform 1 0 2544 0 -1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_79
timestamp 1681708930
transform -1 0 2576 0 -1 570
box -8 -3 32 105
use FILL  FILL_1369
timestamp 1681708930
transform 1 0 2576 0 -1 570
box -8 -3 16 105
use FILL  FILL_1370
timestamp 1681708930
transform 1 0 2584 0 -1 570
box -8 -3 16 105
use XNOR2X1  XNOR2X1_51
timestamp 1681708930
transform -1 0 2648 0 -1 570
box -8 -3 64 105
use FILL  FILL_1371
timestamp 1681708930
transform 1 0 2648 0 -1 570
box -8 -3 16 105
use FILL  FILL_1373
timestamp 1681708930
transform 1 0 2656 0 -1 570
box -8 -3 16 105
use top_mod_new_VIA0  top_mod_new_VIA0_43
timestamp 1681708930
transform 1 0 2712 0 1 470
box -10 -3 10 3
use M3_M2  M3_M2_3443
timestamp 1681708930
transform 1 0 68 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_3444
timestamp 1681708930
transform 1 0 172 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3504
timestamp 1681708930
transform 1 0 188 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3538
timestamp 1681708930
transform 1 0 68 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3539
timestamp 1681708930
transform 1 0 132 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3605
timestamp 1681708930
transform 1 0 156 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3606
timestamp 1681708930
transform 1 0 172 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3607
timestamp 1681708930
transform 1 0 188 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3513
timestamp 1681708930
transform 1 0 132 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3514
timestamp 1681708930
transform 1 0 188 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3445
timestamp 1681708930
transform 1 0 220 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3540
timestamp 1681708930
transform 1 0 220 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3541
timestamp 1681708930
transform 1 0 228 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3542
timestamp 1681708930
transform 1 0 284 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3468
timestamp 1681708930
transform 1 0 308 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3417
timestamp 1681708930
transform 1 0 348 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_3505
timestamp 1681708930
transform 1 0 348 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_3446
timestamp 1681708930
transform 1 0 356 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3506
timestamp 1681708930
transform 1 0 380 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3543
timestamp 1681708930
transform 1 0 332 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3608
timestamp 1681708930
transform 1 0 220 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3609
timestamp 1681708930
transform 1 0 308 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3610
timestamp 1681708930
transform 1 0 324 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3515
timestamp 1681708930
transform 1 0 220 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3516
timestamp 1681708930
transform 1 0 236 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3517
timestamp 1681708930
transform 1 0 284 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3495
timestamp 1681708930
transform 1 0 332 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_3447
timestamp 1681708930
transform 1 0 396 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3544
timestamp 1681708930
transform 1 0 364 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3545
timestamp 1681708930
transform 1 0 380 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3546
timestamp 1681708930
transform 1 0 444 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3611
timestamp 1681708930
transform 1 0 348 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3612
timestamp 1681708930
transform 1 0 356 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3496
timestamp 1681708930
transform 1 0 364 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_3469
timestamp 1681708930
transform 1 0 468 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3418
timestamp 1681708930
transform 1 0 580 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3448
timestamp 1681708930
transform 1 0 564 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3547
timestamp 1681708930
transform 1 0 484 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3548
timestamp 1681708930
transform 1 0 500 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3549
timestamp 1681708930
transform 1 0 516 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3550
timestamp 1681708930
transform 1 0 524 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3551
timestamp 1681708930
transform 1 0 540 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3613
timestamp 1681708930
transform 1 0 380 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3614
timestamp 1681708930
transform 1 0 468 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3518
timestamp 1681708930
transform 1 0 348 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3528
timestamp 1681708930
transform 1 0 340 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3529
timestamp 1681708930
transform 1 0 380 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3470
timestamp 1681708930
transform 1 0 548 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_3552
timestamp 1681708930
transform 1 0 556 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3553
timestamp 1681708930
transform 1 0 580 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3554
timestamp 1681708930
transform 1 0 604 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3615
timestamp 1681708930
transform 1 0 492 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3616
timestamp 1681708930
transform 1 0 508 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3497
timestamp 1681708930
transform 1 0 524 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_3617
timestamp 1681708930
transform 1 0 532 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3618
timestamp 1681708930
transform 1 0 548 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3619
timestamp 1681708930
transform 1 0 564 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3620
timestamp 1681708930
transform 1 0 572 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3621
timestamp 1681708930
transform 1 0 588 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3622
timestamp 1681708930
transform 1 0 596 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3519
timestamp 1681708930
transform 1 0 516 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3530
timestamp 1681708930
transform 1 0 508 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3531
timestamp 1681708930
transform 1 0 548 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3532
timestamp 1681708930
transform 1 0 564 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_3507
timestamp 1681708930
transform 1 0 716 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3555
timestamp 1681708930
transform 1 0 676 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3556
timestamp 1681708930
transform 1 0 708 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3623
timestamp 1681708930
transform 1 0 612 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3624
timestamp 1681708930
transform 1 0 628 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3498
timestamp 1681708930
transform 1 0 676 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_3499
timestamp 1681708930
transform 1 0 708 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_3625
timestamp 1681708930
transform 1 0 716 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3533
timestamp 1681708930
transform 1 0 668 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3449
timestamp 1681708930
transform 1 0 740 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_3400
timestamp 1681708930
transform 1 0 860 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_3409
timestamp 1681708930
transform 1 0 844 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3450
timestamp 1681708930
transform 1 0 844 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3557
timestamp 1681708930
transform 1 0 740 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3558
timestamp 1681708930
transform 1 0 748 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3559
timestamp 1681708930
transform 1 0 804 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3471
timestamp 1681708930
transform 1 0 828 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3401
timestamp 1681708930
transform 1 0 932 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_3410
timestamp 1681708930
transform 1 0 916 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3419
timestamp 1681708930
transform 1 0 900 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_3508
timestamp 1681708930
transform 1 0 868 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_3451
timestamp 1681708930
transform 1 0 876 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3509
timestamp 1681708930
transform 1 0 900 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3560
timestamp 1681708930
transform 1 0 852 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3472
timestamp 1681708930
transform 1 0 860 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_3626
timestamp 1681708930
transform 1 0 740 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3627
timestamp 1681708930
transform 1 0 828 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3628
timestamp 1681708930
transform 1 0 844 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3534
timestamp 1681708930
transform 1 0 804 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3500
timestamp 1681708930
transform 1 0 852 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_3561
timestamp 1681708930
transform 1 0 884 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3629
timestamp 1681708930
transform 1 0 868 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3630
timestamp 1681708930
transform 1 0 876 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3501
timestamp 1681708930
transform 1 0 884 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_3452
timestamp 1681708930
transform 1 0 924 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3562
timestamp 1681708930
transform 1 0 908 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3473
timestamp 1681708930
transform 1 0 916 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_3563
timestamp 1681708930
transform 1 0 924 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3631
timestamp 1681708930
transform 1 0 900 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3632
timestamp 1681708930
transform 1 0 916 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3633
timestamp 1681708930
transform 1 0 932 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3535
timestamp 1681708930
transform 1 0 868 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_3564
timestamp 1681708930
transform 1 0 964 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3502
timestamp 1681708930
transform 1 0 964 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_3411
timestamp 1681708930
transform 1 0 980 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3420
timestamp 1681708930
transform 1 0 996 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3453
timestamp 1681708930
transform 1 0 980 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3565
timestamp 1681708930
transform 1 0 972 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3566
timestamp 1681708930
transform 1 0 996 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3474
timestamp 1681708930
transform 1 0 1004 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_3567
timestamp 1681708930
transform 1 0 1012 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3568
timestamp 1681708930
transform 1 0 1020 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3634
timestamp 1681708930
transform 1 0 988 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3635
timestamp 1681708930
transform 1 0 1004 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3536
timestamp 1681708930
transform 1 0 988 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3402
timestamp 1681708930
transform 1 0 1044 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_3454
timestamp 1681708930
transform 1 0 1044 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3636
timestamp 1681708930
transform 1 0 1028 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3537
timestamp 1681708930
transform 1 0 1052 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3412
timestamp 1681708930
transform 1 0 1084 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_3510
timestamp 1681708930
transform 1 0 1084 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3637
timestamp 1681708930
transform 1 0 1100 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3538
timestamp 1681708930
transform 1 0 1100 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_3492
timestamp 1681708930
transform 1 0 1116 0 1 435
box -2 -2 2 2
use M3_M2  M3_M2_3455
timestamp 1681708930
transform 1 0 1116 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3511
timestamp 1681708930
transform 1 0 1132 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3569
timestamp 1681708930
transform 1 0 1124 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3570
timestamp 1681708930
transform 1 0 1140 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3503
timestamp 1681708930
transform 1 0 1116 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_3520
timestamp 1681708930
transform 1 0 1132 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3404
timestamp 1681708930
transform 1 0 1164 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_3475
timestamp 1681708930
transform 1 0 1164 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3421
timestamp 1681708930
transform 1 0 1188 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_3512
timestamp 1681708930
transform 1 0 1188 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3638
timestamp 1681708930
transform 1 0 1164 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3639
timestamp 1681708930
transform 1 0 1172 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3504
timestamp 1681708930
transform 1 0 1180 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_3675
timestamp 1681708930
transform 1 0 1180 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_3539
timestamp 1681708930
transform 1 0 1172 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3405
timestamp 1681708930
transform 1 0 1220 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_3413
timestamp 1681708930
transform 1 0 1228 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3456
timestamp 1681708930
transform 1 0 1236 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3571
timestamp 1681708930
transform 1 0 1204 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3572
timestamp 1681708930
transform 1 0 1220 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3573
timestamp 1681708930
transform 1 0 1236 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3505
timestamp 1681708930
transform 1 0 1204 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_3406
timestamp 1681708930
transform 1 0 1292 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_3414
timestamp 1681708930
transform 1 0 1276 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3422
timestamp 1681708930
transform 1 0 1284 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_3574
timestamp 1681708930
transform 1 0 1260 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3640
timestamp 1681708930
transform 1 0 1212 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3641
timestamp 1681708930
transform 1 0 1228 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3642
timestamp 1681708930
transform 1 0 1252 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3476
timestamp 1681708930
transform 1 0 1268 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_3575
timestamp 1681708930
transform 1 0 1284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3643
timestamp 1681708930
transform 1 0 1268 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3644
timestamp 1681708930
transform 1 0 1292 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3513
timestamp 1681708930
transform 1 0 1308 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3576
timestamp 1681708930
transform 1 0 1316 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3423
timestamp 1681708930
transform 1 0 1356 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_3493
timestamp 1681708930
transform 1 0 1364 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_3514
timestamp 1681708930
transform 1 0 1364 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3577
timestamp 1681708930
transform 1 0 1356 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3477
timestamp 1681708930
transform 1 0 1364 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_3578
timestamp 1681708930
transform 1 0 1372 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3506
timestamp 1681708930
transform 1 0 1372 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_3478
timestamp 1681708930
transform 1 0 1388 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_3645
timestamp 1681708930
transform 1 0 1380 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3646
timestamp 1681708930
transform 1 0 1388 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3540
timestamp 1681708930
transform 1 0 1348 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3507
timestamp 1681708930
transform 1 0 1396 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_3515
timestamp 1681708930
transform 1 0 1420 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_3424
timestamp 1681708930
transform 1 0 1452 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_3494
timestamp 1681708930
transform 1 0 1460 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_3516
timestamp 1681708930
transform 1 0 1452 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3579
timestamp 1681708930
transform 1 0 1436 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3425
timestamp 1681708930
transform 1 0 1476 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_3517
timestamp 1681708930
transform 1 0 1476 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3580
timestamp 1681708930
transform 1 0 1468 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3647
timestamp 1681708930
transform 1 0 1444 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3521
timestamp 1681708930
transform 1 0 1436 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_3648
timestamp 1681708930
transform 1 0 1484 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3676
timestamp 1681708930
transform 1 0 1484 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_3426
timestamp 1681708930
transform 1 0 1524 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3457
timestamp 1681708930
transform 1 0 1508 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3581
timestamp 1681708930
transform 1 0 1508 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3649
timestamp 1681708930
transform 1 0 1500 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3522
timestamp 1681708930
transform 1 0 1500 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3458
timestamp 1681708930
transform 1 0 1556 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3582
timestamp 1681708930
transform 1 0 1564 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3650
timestamp 1681708930
transform 1 0 1556 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3479
timestamp 1681708930
transform 1 0 1572 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3427
timestamp 1681708930
transform 1 0 1588 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_3495
timestamp 1681708930
transform 1 0 1604 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_3496
timestamp 1681708930
transform 1 0 1612 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_3518
timestamp 1681708930
transform 1 0 1588 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3519
timestamp 1681708930
transform 1 0 1596 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3583
timestamp 1681708930
transform 1 0 1580 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3651
timestamp 1681708930
transform 1 0 1572 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3523
timestamp 1681708930
transform 1 0 1572 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3459
timestamp 1681708930
transform 1 0 1604 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3520
timestamp 1681708930
transform 1 0 1620 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3584
timestamp 1681708930
transform 1 0 1604 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3480
timestamp 1681708930
transform 1 0 1612 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3428
timestamp 1681708930
transform 1 0 1652 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_3585
timestamp 1681708930
transform 1 0 1644 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3481
timestamp 1681708930
transform 1 0 1660 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_3652
timestamp 1681708930
transform 1 0 1676 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3429
timestamp 1681708930
transform 1 0 1788 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3460
timestamp 1681708930
transform 1 0 1764 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_3461
timestamp 1681708930
transform 1 0 1780 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3497
timestamp 1681708930
transform 1 0 1860 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_3521
timestamp 1681708930
transform 1 0 1844 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3586
timestamp 1681708930
transform 1 0 1780 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3587
timestamp 1681708930
transform 1 0 1788 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3482
timestamp 1681708930
transform 1 0 1812 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3508
timestamp 1681708930
transform 1 0 1780 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_3653
timestamp 1681708930
transform 1 0 1788 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3524
timestamp 1681708930
transform 1 0 1780 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_3654
timestamp 1681708930
transform 1 0 1836 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3525
timestamp 1681708930
transform 1 0 1836 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3541
timestamp 1681708930
transform 1 0 1844 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3430
timestamp 1681708930
transform 1 0 1868 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_3522
timestamp 1681708930
transform 1 0 1868 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3588
timestamp 1681708930
transform 1 0 1884 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3542
timestamp 1681708930
transform 1 0 1876 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_3655
timestamp 1681708930
transform 1 0 1892 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3656
timestamp 1681708930
transform 1 0 1900 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3543
timestamp 1681708930
transform 1 0 1900 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3403
timestamp 1681708930
transform 1 0 1980 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_3431
timestamp 1681708930
transform 1 0 1964 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_3498
timestamp 1681708930
transform 1 0 1972 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_3523
timestamp 1681708930
transform 1 0 1956 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3524
timestamp 1681708930
transform 1 0 1980 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_3432
timestamp 1681708930
transform 1 0 2020 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_3589
timestamp 1681708930
transform 1 0 1964 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3590
timestamp 1681708930
transform 1 0 1988 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3657
timestamp 1681708930
transform 1 0 1948 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3483
timestamp 1681708930
transform 1 0 2004 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_3591
timestamp 1681708930
transform 1 0 2020 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3658
timestamp 1681708930
transform 1 0 2004 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3677
timestamp 1681708930
transform 1 0 1988 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_3499
timestamp 1681708930
transform 1 0 2052 0 1 435
box -2 -2 2 2
use M3_M2  M3_M2_3433
timestamp 1681708930
transform 1 0 2060 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_3525
timestamp 1681708930
transform 1 0 2044 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_3434
timestamp 1681708930
transform 1 0 2084 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3435
timestamp 1681708930
transform 1 0 2132 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_3526
timestamp 1681708930
transform 1 0 2068 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_3462
timestamp 1681708930
transform 1 0 2108 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_3463
timestamp 1681708930
transform 1 0 2124 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3592
timestamp 1681708930
transform 1 0 2060 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3678
timestamp 1681708930
transform 1 0 2036 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_3484
timestamp 1681708930
transform 1 0 2068 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_3593
timestamp 1681708930
transform 1 0 2100 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3594
timestamp 1681708930
transform 1 0 2108 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3659
timestamp 1681708930
transform 1 0 2076 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3544
timestamp 1681708930
transform 1 0 2060 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3436
timestamp 1681708930
transform 1 0 2212 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3437
timestamp 1681708930
transform 1 0 2244 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3485
timestamp 1681708930
transform 1 0 2148 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3486
timestamp 1681708930
transform 1 0 2180 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_3595
timestamp 1681708930
transform 1 0 2212 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3660
timestamp 1681708930
transform 1 0 2124 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3661
timestamp 1681708930
transform 1 0 2132 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3526
timestamp 1681708930
transform 1 0 2132 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3545
timestamp 1681708930
transform 1 0 2084 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3546
timestamp 1681708930
transform 1 0 2124 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_3662
timestamp 1681708930
transform 1 0 2180 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3663
timestamp 1681708930
transform 1 0 2188 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3487
timestamp 1681708930
transform 1 0 2244 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_3500
timestamp 1681708930
transform 1 0 2316 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_3527
timestamp 1681708930
transform 1 0 2300 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3596
timestamp 1681708930
transform 1 0 2268 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3664
timestamp 1681708930
transform 1 0 2236 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3665
timestamp 1681708930
transform 1 0 2244 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3527
timestamp 1681708930
transform 1 0 2236 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3488
timestamp 1681708930
transform 1 0 2292 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_3528
timestamp 1681708930
transform 1 0 2324 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3597
timestamp 1681708930
transform 1 0 2308 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3666
timestamp 1681708930
transform 1 0 2292 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3547
timestamp 1681708930
transform 1 0 2292 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3489
timestamp 1681708930
transform 1 0 2324 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_3598
timestamp 1681708930
transform 1 0 2332 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3509
timestamp 1681708930
transform 1 0 2332 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_3548
timestamp 1681708930
transform 1 0 2340 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3464
timestamp 1681708930
transform 1 0 2380 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3529
timestamp 1681708930
transform 1 0 2388 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3667
timestamp 1681708930
transform 1 0 2372 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3679
timestamp 1681708930
transform 1 0 2388 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_3415
timestamp 1681708930
transform 1 0 2412 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_3501
timestamp 1681708930
transform 1 0 2412 0 1 435
box -2 -2 2 2
use M3_M2  M3_M2_3438
timestamp 1681708930
transform 1 0 2428 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_3502
timestamp 1681708930
transform 1 0 2436 0 1 435
box -2 -2 2 2
use M3_M2  M3_M2_3465
timestamp 1681708930
transform 1 0 2404 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3530
timestamp 1681708930
transform 1 0 2412 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3531
timestamp 1681708930
transform 1 0 2428 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3599
timestamp 1681708930
transform 1 0 2412 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3549
timestamp 1681708930
transform 1 0 2404 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3466
timestamp 1681708930
transform 1 0 2444 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_3532
timestamp 1681708930
transform 1 0 2452 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3533
timestamp 1681708930
transform 1 0 2460 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3600
timestamp 1681708930
transform 1 0 2444 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3467
timestamp 1681708930
transform 1 0 2476 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_3439
timestamp 1681708930
transform 1 0 2500 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3490
timestamp 1681708930
transform 1 0 2468 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3491
timestamp 1681708930
transform 1 0 2484 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_3601
timestamp 1681708930
transform 1 0 2500 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3492
timestamp 1681708930
transform 1 0 2508 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_3668
timestamp 1681708930
transform 1 0 2460 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3669
timestamp 1681708930
transform 1 0 2484 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3670
timestamp 1681708930
transform 1 0 2492 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3510
timestamp 1681708930
transform 1 0 2500 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_3671
timestamp 1681708930
transform 1 0 2508 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3680
timestamp 1681708930
transform 1 0 2508 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_3407
timestamp 1681708930
transform 1 0 2556 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_3416
timestamp 1681708930
transform 1 0 2572 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3440
timestamp 1681708930
transform 1 0 2564 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_3503
timestamp 1681708930
transform 1 0 2580 0 1 435
box -2 -2 2 2
use M3_M2  M3_M2_3441
timestamp 1681708930
transform 1 0 2588 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3442
timestamp 1681708930
transform 1 0 2604 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_3534
timestamp 1681708930
transform 1 0 2556 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3535
timestamp 1681708930
transform 1 0 2564 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3536
timestamp 1681708930
transform 1 0 2588 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3602
timestamp 1681708930
transform 1 0 2540 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3493
timestamp 1681708930
transform 1 0 2548 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_3603
timestamp 1681708930
transform 1 0 2556 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3494
timestamp 1681708930
transform 1 0 2564 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_3604
timestamp 1681708930
transform 1 0 2572 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_3511
timestamp 1681708930
transform 1 0 2540 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_3672
timestamp 1681708930
transform 1 0 2596 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_3408
timestamp 1681708930
transform 1 0 2628 0 1 455
box -3 -3 3 3
use M2_M1  M2_M1_3673
timestamp 1681708930
transform 1 0 2620 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3674
timestamp 1681708930
transform 1 0 2628 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3537
timestamp 1681708930
transform 1 0 2652 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_3512
timestamp 1681708930
transform 1 0 2652 0 1 405
box -3 -3 3 3
use top_mod_new_VIA0  top_mod_new_VIA0_44
timestamp 1681708930
transform 1 0 48 0 1 370
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_86
timestamp 1681708930
transform -1 0 168 0 1 370
box -8 -3 104 105
use NAND2X1  NAND2X1_82
timestamp 1681708930
transform 1 0 168 0 1 370
box -8 -3 32 105
use OAI21X1  OAI21X1_88
timestamp 1681708930
transform -1 0 224 0 1 370
box -8 -3 34 105
use M3_M2  M3_M2_3550
timestamp 1681708930
transform 1 0 308 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_88
timestamp 1681708930
transform -1 0 320 0 1 370
box -8 -3 104 105
use M3_M2  M3_M2_3551
timestamp 1681708930
transform 1 0 340 0 1 375
box -3 -3 3 3
use OAI21X1  OAI21X1_89
timestamp 1681708930
transform 1 0 320 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_90
timestamp 1681708930
transform 1 0 352 0 1 370
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_89
timestamp 1681708930
transform -1 0 480 0 1 370
box -8 -3 104 105
use AOI22X1  AOI22X1_87
timestamp 1681708930
transform 1 0 480 0 1 370
box -8 -3 46 105
use M3_M2  M3_M2_3552
timestamp 1681708930
transform 1 0 556 0 1 375
box -3 -3 3 3
use AOI22X1  AOI22X1_88
timestamp 1681708930
transform 1 0 520 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_89
timestamp 1681708930
transform 1 0 560 0 1 370
box -8 -3 46 105
use INVX2  INVX2_232
timestamp 1681708930
transform -1 0 616 0 1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_90
timestamp 1681708930
transform 1 0 616 0 1 370
box -8 -3 104 105
use OAI21X1  OAI21X1_91
timestamp 1681708930
transform -1 0 744 0 1 370
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_91
timestamp 1681708930
transform -1 0 840 0 1 370
box -8 -3 104 105
use OAI21X1  OAI21X1_92
timestamp 1681708930
transform 1 0 840 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_93
timestamp 1681708930
transform 1 0 872 0 1 370
box -8 -3 34 105
use AOI22X1  AOI22X1_90
timestamp 1681708930
transform 1 0 904 0 1 370
box -8 -3 46 105
use FILL  FILL_1374
timestamp 1681708930
transform 1 0 944 0 1 370
box -8 -3 16 105
use FILL  FILL_1375
timestamp 1681708930
transform 1 0 952 0 1 370
box -8 -3 16 105
use FILL  FILL_1407
timestamp 1681708930
transform 1 0 960 0 1 370
box -8 -3 16 105
use FILL  FILL_1409
timestamp 1681708930
transform 1 0 968 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_92
timestamp 1681708930
transform -1 0 1016 0 1 370
box -8 -3 46 105
use M3_M2  M3_M2_3553
timestamp 1681708930
transform 1 0 1028 0 1 375
box -3 -3 3 3
use FILL  FILL_1410
timestamp 1681708930
transform 1 0 1016 0 1 370
box -8 -3 16 105
use XOR2X1  XOR2X1_187
timestamp 1681708930
transform -1 0 1080 0 1 370
box -8 -3 64 105
use FILL  FILL_1411
timestamp 1681708930
transform 1 0 1080 0 1 370
box -8 -3 16 105
use FILL  FILL_1412
timestamp 1681708930
transform 1 0 1088 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_3554
timestamp 1681708930
transform 1 0 1108 0 1 375
box -3 -3 3 3
use FILL  FILL_1413
timestamp 1681708930
transform 1 0 1096 0 1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_128
timestamp 1681708930
transform -1 0 1136 0 1 370
box -8 -3 40 105
use OR2X1  OR2X1_23
timestamp 1681708930
transform -1 0 1168 0 1 370
box -8 -3 40 105
use FILL  FILL_1414
timestamp 1681708930
transform 1 0 1168 0 1 370
box -8 -3 16 105
use FILL  FILL_1415
timestamp 1681708930
transform 1 0 1176 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_98
timestamp 1681708930
transform -1 0 1216 0 1 370
box -8 -3 34 105
use AOI22X1  AOI22X1_93
timestamp 1681708930
transform 1 0 1216 0 1 370
box -8 -3 46 105
use FILL  FILL_1416
timestamp 1681708930
transform 1 0 1256 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_94
timestamp 1681708930
transform -1 0 1304 0 1 370
box -8 -3 46 105
use FILL  FILL_1417
timestamp 1681708930
transform 1 0 1304 0 1 370
box -8 -3 16 105
use FILL  FILL_1418
timestamp 1681708930
transform 1 0 1312 0 1 370
box -8 -3 16 105
use FILL  FILL_1419
timestamp 1681708930
transform 1 0 1320 0 1 370
box -8 -3 16 105
use FILL  FILL_1432
timestamp 1681708930
transform 1 0 1328 0 1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_129
timestamp 1681708930
transform -1 0 1368 0 1 370
box -8 -3 40 105
use INVX2  INVX2_238
timestamp 1681708930
transform -1 0 1384 0 1 370
box -9 -3 26 105
use FILL  FILL_1433
timestamp 1681708930
transform 1 0 1384 0 1 370
box -8 -3 16 105
use FILL  FILL_1434
timestamp 1681708930
transform 1 0 1392 0 1 370
box -8 -3 16 105
use FILL  FILL_1435
timestamp 1681708930
transform 1 0 1400 0 1 370
box -8 -3 16 105
use FILL  FILL_1436
timestamp 1681708930
transform 1 0 1408 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_99
timestamp 1681708930
transform -1 0 1448 0 1 370
box -8 -3 34 105
use NAND3X1  NAND3X1_130
timestamp 1681708930
transform -1 0 1480 0 1 370
box -8 -3 40 105
use NOR2X1  NOR2X1_80
timestamp 1681708930
transform 1 0 1480 0 1 370
box -8 -3 32 105
use XNOR2X1  XNOR2X1_52
timestamp 1681708930
transform 1 0 1504 0 1 370
box -8 -3 64 105
use FILL  FILL_1437
timestamp 1681708930
transform 1 0 1560 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_85
timestamp 1681708930
transform 1 0 1568 0 1 370
box -8 -3 32 105
use NAND3X1  NAND3X1_131
timestamp 1681708930
transform 1 0 1592 0 1 370
box -8 -3 40 105
use FILL  FILL_1438
timestamp 1681708930
transform 1 0 1624 0 1 370
box -8 -3 16 105
use FILL  FILL_1439
timestamp 1681708930
transform 1 0 1632 0 1 370
box -8 -3 16 105
use FILL  FILL_1440
timestamp 1681708930
transform 1 0 1640 0 1 370
box -8 -3 16 105
use FILL  FILL_1441
timestamp 1681708930
transform 1 0 1648 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_3555
timestamp 1681708930
transform 1 0 1668 0 1 375
box -3 -3 3 3
use FILL  FILL_1442
timestamp 1681708930
transform 1 0 1656 0 1 370
box -8 -3 16 105
use FILL  FILL_1443
timestamp 1681708930
transform 1 0 1664 0 1 370
box -8 -3 16 105
use FILL  FILL_1444
timestamp 1681708930
transform 1 0 1672 0 1 370
box -8 -3 16 105
use FILL  FILL_1445
timestamp 1681708930
transform 1 0 1680 0 1 370
box -8 -3 16 105
use FILL  FILL_1446
timestamp 1681708930
transform 1 0 1688 0 1 370
box -8 -3 16 105
use FILL  FILL_1447
timestamp 1681708930
transform 1 0 1696 0 1 370
box -8 -3 16 105
use FILL  FILL_1448
timestamp 1681708930
transform 1 0 1704 0 1 370
box -8 -3 16 105
use FILL  FILL_1449
timestamp 1681708930
transform 1 0 1712 0 1 370
box -8 -3 16 105
use FILL  FILL_1450
timestamp 1681708930
transform 1 0 1720 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_3556
timestamp 1681708930
transform 1 0 1772 0 1 375
box -3 -3 3 3
use XOR2X1  XOR2X1_192
timestamp 1681708930
transform -1 0 1784 0 1 370
box -8 -3 64 105
use M3_M2  M3_M2_3557
timestamp 1681708930
transform 1 0 1812 0 1 375
box -3 -3 3 3
use XOR2X1  XOR2X1_193
timestamp 1681708930
transform -1 0 1840 0 1 370
box -8 -3 64 105
use NAND3X1  NAND3X1_132
timestamp 1681708930
transform -1 0 1872 0 1 370
box -8 -3 40 105
use INVX2  INVX2_239
timestamp 1681708930
transform -1 0 1888 0 1 370
box -9 -3 26 105
use FILL  FILL_1451
timestamp 1681708930
transform 1 0 1888 0 1 370
box -8 -3 16 105
use XOR2X1  XOR2X1_194
timestamp 1681708930
transform -1 0 1952 0 1 370
box -8 -3 64 105
use NAND3X1  NAND3X1_133
timestamp 1681708930
transform 1 0 1952 0 1 370
box -8 -3 40 105
use AOI21X1  AOI21X1_49
timestamp 1681708930
transform -1 0 2016 0 1 370
box -7 -3 39 105
use NOR2X1  NOR2X1_81
timestamp 1681708930
transform -1 0 2040 0 1 370
box -8 -3 32 105
use M3_M2  M3_M2_3558
timestamp 1681708930
transform 1 0 2052 0 1 375
box -3 -3 3 3
use NAND3X1  NAND3X1_134
timestamp 1681708930
transform -1 0 2072 0 1 370
box -8 -3 40 105
use XOR2X1  XOR2X1_195
timestamp 1681708930
transform 1 0 2072 0 1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_196
timestamp 1681708930
transform -1 0 2184 0 1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_197
timestamp 1681708930
transform 1 0 2184 0 1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_198
timestamp 1681708930
transform 1 0 2240 0 1 370
box -8 -3 64 105
use NAND3X1  NAND3X1_135
timestamp 1681708930
transform 1 0 2296 0 1 370
box -8 -3 40 105
use FILL  FILL_1452
timestamp 1681708930
transform 1 0 2328 0 1 370
box -8 -3 16 105
use FILL  FILL_1453
timestamp 1681708930
transform 1 0 2336 0 1 370
box -8 -3 16 105
use FILL  FILL_1484
timestamp 1681708930
transform 1 0 2344 0 1 370
box -8 -3 16 105
use OR2X1  OR2X1_26
timestamp 1681708930
transform -1 0 2384 0 1 370
box -8 -3 40 105
use FILL  FILL_1485
timestamp 1681708930
transform 1 0 2384 0 1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_141
timestamp 1681708930
transform -1 0 2424 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_142
timestamp 1681708930
transform -1 0 2456 0 1 370
box -8 -3 40 105
use OAI21X1  OAI21X1_105
timestamp 1681708930
transform -1 0 2488 0 1 370
box -8 -3 34 105
use INVX2  INVX2_244
timestamp 1681708930
transform 1 0 2488 0 1 370
box -9 -3 26 105
use NOR2X1  NOR2X1_84
timestamp 1681708930
transform 1 0 2504 0 1 370
box -8 -3 32 105
use FILL  FILL_1486
timestamp 1681708930
transform 1 0 2528 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_88
timestamp 1681708930
transform 1 0 2536 0 1 370
box -8 -3 32 105
use NAND3X1  NAND3X1_143
timestamp 1681708930
transform 1 0 2560 0 1 370
box -8 -3 40 105
use OAI21X1  OAI21X1_106
timestamp 1681708930
transform -1 0 2624 0 1 370
box -8 -3 34 105
use FILL  FILL_1487
timestamp 1681708930
transform 1 0 2624 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_89
timestamp 1681708930
transform 1 0 2632 0 1 370
box -8 -3 32 105
use FILL  FILL_1488
timestamp 1681708930
transform 1 0 2656 0 1 370
box -8 -3 16 105
use top_mod_new_VIA0  top_mod_new_VIA0_45
timestamp 1681708930
transform 1 0 2688 0 1 370
box -10 -3 10 3
use M3_M2  M3_M2_3593
timestamp 1681708930
transform 1 0 132 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3617
timestamp 1681708930
transform 1 0 68 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3594
timestamp 1681708930
transform 1 0 188 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_3690
timestamp 1681708930
transform 1 0 156 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3691
timestamp 1681708930
transform 1 0 172 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3761
timestamp 1681708930
transform 1 0 68 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3762
timestamp 1681708930
transform 1 0 132 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3618
timestamp 1681708930
transform 1 0 180 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_3692
timestamp 1681708930
transform 1 0 188 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3822
timestamp 1681708930
transform 1 0 188 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_3559
timestamp 1681708930
transform 1 0 228 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_3693
timestamp 1681708930
transform 1 0 220 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3694
timestamp 1681708930
transform 1 0 228 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3668
timestamp 1681708930
transform 1 0 220 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3577
timestamp 1681708930
transform 1 0 284 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3619
timestamp 1681708930
transform 1 0 260 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3560
timestamp 1681708930
transform 1 0 308 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_3695
timestamp 1681708930
transform 1 0 300 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3763
timestamp 1681708930
transform 1 0 260 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3764
timestamp 1681708930
transform 1 0 268 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3765
timestamp 1681708930
transform 1 0 284 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3685
timestamp 1681708930
transform 1 0 276 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_3578
timestamp 1681708930
transform 1 0 332 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3595
timestamp 1681708930
transform 1 0 324 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_3696
timestamp 1681708930
transform 1 0 308 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3620
timestamp 1681708930
transform 1 0 316 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_3766
timestamp 1681708930
transform 1 0 316 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3823
timestamp 1681708930
transform 1 0 308 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3767
timestamp 1681708930
transform 1 0 332 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3669
timestamp 1681708930
transform 1 0 332 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_3697
timestamp 1681708930
transform 1 0 372 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3698
timestamp 1681708930
transform 1 0 412 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3579
timestamp 1681708930
transform 1 0 436 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_3699
timestamp 1681708930
transform 1 0 428 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3768
timestamp 1681708930
transform 1 0 420 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3769
timestamp 1681708930
transform 1 0 436 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3670
timestamp 1681708930
transform 1 0 428 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3686
timestamp 1681708930
transform 1 0 428 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_3700
timestamp 1681708930
transform 1 0 460 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3701
timestamp 1681708930
transform 1 0 492 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3824
timestamp 1681708930
transform 1 0 500 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_3561
timestamp 1681708930
transform 1 0 532 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3562
timestamp 1681708930
transform 1 0 572 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3563
timestamp 1681708930
transform 1 0 596 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3596
timestamp 1681708930
transform 1 0 540 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_3702
timestamp 1681708930
transform 1 0 532 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3703
timestamp 1681708930
transform 1 0 556 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3770
timestamp 1681708930
transform 1 0 524 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3580
timestamp 1681708930
transform 1 0 628 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3597
timestamp 1681708930
transform 1 0 580 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3598
timestamp 1681708930
transform 1 0 628 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_3704
timestamp 1681708930
transform 1 0 580 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3599
timestamp 1681708930
transform 1 0 684 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_3705
timestamp 1681708930
transform 1 0 684 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3771
timestamp 1681708930
transform 1 0 548 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3772
timestamp 1681708930
transform 1 0 564 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3773
timestamp 1681708930
transform 1 0 628 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3774
timestamp 1681708930
transform 1 0 668 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3698
timestamp 1681708930
transform 1 0 644 0 1 285
box -3 -3 3 3
use M2_M1  M2_M1_3825
timestamp 1681708930
transform 1 0 684 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_3621
timestamp 1681708930
transform 1 0 716 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_3775
timestamp 1681708930
transform 1 0 716 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3699
timestamp 1681708930
transform 1 0 700 0 1 285
box -3 -3 3 3
use M2_M1  M2_M1_3706
timestamp 1681708930
transform 1 0 740 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3634
timestamp 1681708930
transform 1 0 732 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3581
timestamp 1681708930
transform 1 0 788 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3582
timestamp 1681708930
transform 1 0 884 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3583
timestamp 1681708930
transform 1 0 900 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3600
timestamp 1681708930
transform 1 0 844 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3601
timestamp 1681708930
transform 1 0 892 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_3707
timestamp 1681708930
transform 1 0 796 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3622
timestamp 1681708930
transform 1 0 876 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3623
timestamp 1681708930
transform 1 0 892 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_3708
timestamp 1681708930
transform 1 0 900 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3776
timestamp 1681708930
transform 1 0 844 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3651
timestamp 1681708930
transform 1 0 860 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_3777
timestamp 1681708930
transform 1 0 892 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3778
timestamp 1681708930
transform 1 0 900 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3584
timestamp 1681708930
transform 1 0 964 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3687
timestamp 1681708930
transform 1 0 964 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_3709
timestamp 1681708930
transform 1 0 980 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3710
timestamp 1681708930
transform 1 0 1012 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3564
timestamp 1681708930
transform 1 0 1060 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_3711
timestamp 1681708930
transform 1 0 1052 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3712
timestamp 1681708930
transform 1 0 1060 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3779
timestamp 1681708930
transform 1 0 1028 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3635
timestamp 1681708930
transform 1 0 1036 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_3780
timestamp 1681708930
transform 1 0 1044 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3602
timestamp 1681708930
transform 1 0 1116 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_3713
timestamp 1681708930
transform 1 0 1116 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3714
timestamp 1681708930
transform 1 0 1124 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3781
timestamp 1681708930
transform 1 0 1084 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3782
timestamp 1681708930
transform 1 0 1092 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3652
timestamp 1681708930
transform 1 0 1092 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_3715
timestamp 1681708930
transform 1 0 1140 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3783
timestamp 1681708930
transform 1 0 1132 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3636
timestamp 1681708930
transform 1 0 1164 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3653
timestamp 1681708930
transform 1 0 1140 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3603
timestamp 1681708930
transform 1 0 1212 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_3716
timestamp 1681708930
transform 1 0 1204 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3717
timestamp 1681708930
transform 1 0 1212 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3637
timestamp 1681708930
transform 1 0 1196 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3671
timestamp 1681708930
transform 1 0 1204 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3585
timestamp 1681708930
transform 1 0 1268 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3586
timestamp 1681708930
transform 1 0 1308 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_3718
timestamp 1681708930
transform 1 0 1260 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3719
timestamp 1681708930
transform 1 0 1268 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3784
timestamp 1681708930
transform 1 0 1236 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3638
timestamp 1681708930
transform 1 0 1260 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_3785
timestamp 1681708930
transform 1 0 1292 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3672
timestamp 1681708930
transform 1 0 1252 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3688
timestamp 1681708930
transform 1 0 1236 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_3654
timestamp 1681708930
transform 1 0 1292 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3639
timestamp 1681708930
transform 1 0 1324 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_3826
timestamp 1681708930
transform 1 0 1324 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3720
timestamp 1681708930
transform 1 0 1348 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3565
timestamp 1681708930
transform 1 0 1380 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3624
timestamp 1681708930
transform 1 0 1364 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_3786
timestamp 1681708930
transform 1 0 1372 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3827
timestamp 1681708930
transform 1 0 1372 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_3625
timestamp 1681708930
transform 1 0 1412 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_3787
timestamp 1681708930
transform 1 0 1412 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3828
timestamp 1681708930
transform 1 0 1396 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3847
timestamp 1681708930
transform 1 0 1388 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_3673
timestamp 1681708930
transform 1 0 1396 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3689
timestamp 1681708930
transform 1 0 1388 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_3566
timestamp 1681708930
transform 1 0 1428 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_3681
timestamp 1681708930
transform 1 0 1428 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3788
timestamp 1681708930
transform 1 0 1428 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3829
timestamp 1681708930
transform 1 0 1420 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_3690
timestamp 1681708930
transform 1 0 1428 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_3848
timestamp 1681708930
transform 1 0 1468 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_3691
timestamp 1681708930
transform 1 0 1468 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_3721
timestamp 1681708930
transform 1 0 1492 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3789
timestamp 1681708930
transform 1 0 1548 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3626
timestamp 1681708930
transform 1 0 1572 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3567
timestamp 1681708930
transform 1 0 1596 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_3682
timestamp 1681708930
transform 1 0 1604 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3722
timestamp 1681708930
transform 1 0 1596 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3790
timestamp 1681708930
transform 1 0 1580 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3830
timestamp 1681708930
transform 1 0 1564 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_3627
timestamp 1681708930
transform 1 0 1604 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_3723
timestamp 1681708930
transform 1 0 1620 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3791
timestamp 1681708930
transform 1 0 1604 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3640
timestamp 1681708930
transform 1 0 1612 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_3831
timestamp 1681708930
transform 1 0 1612 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_3628
timestamp 1681708930
transform 1 0 1628 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_3683
timestamp 1681708930
transform 1 0 1660 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3724
timestamp 1681708930
transform 1 0 1652 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3629
timestamp 1681708930
transform 1 0 1668 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_3725
timestamp 1681708930
transform 1 0 1676 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3726
timestamp 1681708930
transform 1 0 1684 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3792
timestamp 1681708930
transform 1 0 1652 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3793
timestamp 1681708930
transform 1 0 1660 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3794
timestamp 1681708930
transform 1 0 1684 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3655
timestamp 1681708930
transform 1 0 1652 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3692
timestamp 1681708930
transform 1 0 1660 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_3641
timestamp 1681708930
transform 1 0 1692 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_3727
timestamp 1681708930
transform 1 0 1716 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3728
timestamp 1681708930
transform 1 0 1724 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3568
timestamp 1681708930
transform 1 0 1772 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_3729
timestamp 1681708930
transform 1 0 1772 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3795
timestamp 1681708930
transform 1 0 1708 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3642
timestamp 1681708930
transform 1 0 1716 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3643
timestamp 1681708930
transform 1 0 1748 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_3796
timestamp 1681708930
transform 1 0 1756 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3797
timestamp 1681708930
transform 1 0 1772 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3832
timestamp 1681708930
transform 1 0 1692 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_3656
timestamp 1681708930
transform 1 0 1708 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_3684
timestamp 1681708930
transform 1 0 1820 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3730
timestamp 1681708930
transform 1 0 1812 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3604
timestamp 1681708930
transform 1 0 1828 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_3833
timestamp 1681708930
transform 1 0 1828 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_3569
timestamp 1681708930
transform 1 0 1876 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3605
timestamp 1681708930
transform 1 0 1852 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3606
timestamp 1681708930
transform 1 0 1868 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_3798
timestamp 1681708930
transform 1 0 1860 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3657
timestamp 1681708930
transform 1 0 1860 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_3849
timestamp 1681708930
transform 1 0 1852 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_3570
timestamp 1681708930
transform 1 0 1892 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3644
timestamp 1681708930
transform 1 0 1892 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3571
timestamp 1681708930
transform 1 0 1948 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3572
timestamp 1681708930
transform 1 0 1964 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_3685
timestamp 1681708930
transform 1 0 1948 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3686
timestamp 1681708930
transform 1 0 1972 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3731
timestamp 1681708930
transform 1 0 1932 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3732
timestamp 1681708930
transform 1 0 1956 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3733
timestamp 1681708930
transform 1 0 1964 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3799
timestamp 1681708930
transform 1 0 1908 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3800
timestamp 1681708930
transform 1 0 1924 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3834
timestamp 1681708930
transform 1 0 1892 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_3645
timestamp 1681708930
transform 1 0 1932 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_3801
timestamp 1681708930
transform 1 0 1956 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3674
timestamp 1681708930
transform 1 0 1924 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_3734
timestamp 1681708930
transform 1 0 1988 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3646
timestamp 1681708930
transform 1 0 1972 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_3802
timestamp 1681708930
transform 1 0 1980 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3573
timestamp 1681708930
transform 1 0 2036 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3587
timestamp 1681708930
transform 1 0 2028 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_3687
timestamp 1681708930
transform 1 0 2028 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3735
timestamp 1681708930
transform 1 0 2028 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3803
timestamp 1681708930
transform 1 0 2012 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3835
timestamp 1681708930
transform 1 0 1996 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_3658
timestamp 1681708930
transform 1 0 2004 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3574
timestamp 1681708930
transform 1 0 2068 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3588
timestamp 1681708930
transform 1 0 2060 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_3736
timestamp 1681708930
transform 1 0 2052 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3647
timestamp 1681708930
transform 1 0 2036 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_3804
timestamp 1681708930
transform 1 0 2044 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3648
timestamp 1681708930
transform 1 0 2052 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3607
timestamp 1681708930
transform 1 0 2084 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3608
timestamp 1681708930
transform 1 0 2100 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_3737
timestamp 1681708930
transform 1 0 2076 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3738
timestamp 1681708930
transform 1 0 2084 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3630
timestamp 1681708930
transform 1 0 2092 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3609
timestamp 1681708930
transform 1 0 2132 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_3739
timestamp 1681708930
transform 1 0 2108 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3740
timestamp 1681708930
transform 1 0 2124 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3741
timestamp 1681708930
transform 1 0 2132 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3805
timestamp 1681708930
transform 1 0 2084 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3806
timestamp 1681708930
transform 1 0 2092 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3807
timestamp 1681708930
transform 1 0 2116 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3836
timestamp 1681708930
transform 1 0 2020 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_3659
timestamp 1681708930
transform 1 0 2044 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_3837
timestamp 1681708930
transform 1 0 2052 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_3660
timestamp 1681708930
transform 1 0 2068 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3661
timestamp 1681708930
transform 1 0 2084 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3675
timestamp 1681708930
transform 1 0 2012 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_3850
timestamp 1681708930
transform 1 0 2020 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_3676
timestamp 1681708930
transform 1 0 2028 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3693
timestamp 1681708930
transform 1 0 2020 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_3662
timestamp 1681708930
transform 1 0 2116 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3677
timestamp 1681708930
transform 1 0 2100 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3694
timestamp 1681708930
transform 1 0 2076 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_3808
timestamp 1681708930
transform 1 0 2140 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3688
timestamp 1681708930
transform 1 0 2212 0 1 345
box -2 -2 2 2
use M3_M2  M3_M2_3649
timestamp 1681708930
transform 1 0 2212 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_3838
timestamp 1681708930
transform 1 0 2220 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_3678
timestamp 1681708930
transform 1 0 2220 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3610
timestamp 1681708930
transform 1 0 2244 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_3742
timestamp 1681708930
transform 1 0 2244 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3743
timestamp 1681708930
transform 1 0 2252 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3611
timestamp 1681708930
transform 1 0 2292 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3612
timestamp 1681708930
transform 1 0 2332 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_3744
timestamp 1681708930
transform 1 0 2308 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3631
timestamp 1681708930
transform 1 0 2316 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3575
timestamp 1681708930
transform 1 0 2348 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_3745
timestamp 1681708930
transform 1 0 2332 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3632
timestamp 1681708930
transform 1 0 2340 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_3746
timestamp 1681708930
transform 1 0 2348 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3809
timestamp 1681708930
transform 1 0 2252 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3810
timestamp 1681708930
transform 1 0 2260 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3811
timestamp 1681708930
transform 1 0 2284 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3812
timestamp 1681708930
transform 1 0 2300 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3813
timestamp 1681708930
transform 1 0 2316 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3814
timestamp 1681708930
transform 1 0 2332 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3815
timestamp 1681708930
transform 1 0 2340 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3663
timestamp 1681708930
transform 1 0 2252 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_3839
timestamp 1681708930
transform 1 0 2268 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3840
timestamp 1681708930
transform 1 0 2292 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_3679
timestamp 1681708930
transform 1 0 2268 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3680
timestamp 1681708930
transform 1 0 2284 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3664
timestamp 1681708930
transform 1 0 2316 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3665
timestamp 1681708930
transform 1 0 2332 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_3851
timestamp 1681708930
transform 1 0 2292 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_3695
timestamp 1681708930
transform 1 0 2260 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_3696
timestamp 1681708930
transform 1 0 2284 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_3697
timestamp 1681708930
transform 1 0 2300 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_3700
timestamp 1681708930
transform 1 0 2292 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_3681
timestamp 1681708930
transform 1 0 2332 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3701
timestamp 1681708930
transform 1 0 2332 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_3589
timestamp 1681708930
transform 1 0 2380 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3613
timestamp 1681708930
transform 1 0 2372 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_3689
timestamp 1681708930
transform 1 0 2380 0 1 345
box -2 -2 2 2
use M3_M2  M3_M2_3614
timestamp 1681708930
transform 1 0 2388 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_3816
timestamp 1681708930
transform 1 0 2364 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3702
timestamp 1681708930
transform 1 0 2348 0 1 285
box -3 -3 3 3
use M2_M1  M2_M1_3747
timestamp 1681708930
transform 1 0 2372 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3633
timestamp 1681708930
transform 1 0 2380 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3590
timestamp 1681708930
transform 1 0 2412 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_3748
timestamp 1681708930
transform 1 0 2388 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3749
timestamp 1681708930
transform 1 0 2396 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3750
timestamp 1681708930
transform 1 0 2412 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3666
timestamp 1681708930
transform 1 0 2396 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_3841
timestamp 1681708930
transform 1 0 2404 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_3576
timestamp 1681708930
transform 1 0 2452 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3615
timestamp 1681708930
transform 1 0 2444 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_3751
timestamp 1681708930
transform 1 0 2444 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3752
timestamp 1681708930
transform 1 0 2452 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3817
timestamp 1681708930
transform 1 0 2436 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3842
timestamp 1681708930
transform 1 0 2428 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3852
timestamp 1681708930
transform 1 0 2404 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_3853
timestamp 1681708930
transform 1 0 2420 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_3682
timestamp 1681708930
transform 1 0 2428 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_3753
timestamp 1681708930
transform 1 0 2468 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3754
timestamp 1681708930
transform 1 0 2484 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_3650
timestamp 1681708930
transform 1 0 2484 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3591
timestamp 1681708930
transform 1 0 2532 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_3755
timestamp 1681708930
transform 1 0 2516 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3756
timestamp 1681708930
transform 1 0 2524 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3818
timestamp 1681708930
transform 1 0 2492 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3819
timestamp 1681708930
transform 1 0 2508 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_3667
timestamp 1681708930
transform 1 0 2476 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_3843
timestamp 1681708930
transform 1 0 2484 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3844
timestamp 1681708930
transform 1 0 2492 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_3683
timestamp 1681708930
transform 1 0 2492 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3592
timestamp 1681708930
transform 1 0 2596 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3616
timestamp 1681708930
transform 1 0 2572 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_3757
timestamp 1681708930
transform 1 0 2572 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3758
timestamp 1681708930
transform 1 0 2596 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3759
timestamp 1681708930
transform 1 0 2604 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3760
timestamp 1681708930
transform 1 0 2660 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3820
timestamp 1681708930
transform 1 0 2556 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3845
timestamp 1681708930
transform 1 0 2540 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_3684
timestamp 1681708930
transform 1 0 2548 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_3821
timestamp 1681708930
transform 1 0 2580 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3846
timestamp 1681708930
transform 1 0 2572 0 1 315
box -2 -2 2 2
use top_mod_new_VIA0  top_mod_new_VIA0_46
timestamp 1681708930
transform 1 0 24 0 1 270
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_87
timestamp 1681708930
transform -1 0 168 0 -1 370
box -8 -3 104 105
use NAND2X1  NAND2X1_83
timestamp 1681708930
transform 1 0 168 0 -1 370
box -8 -3 32 105
use OAI21X1  OAI21X1_94
timestamp 1681708930
transform -1 0 224 0 -1 370
box -8 -3 34 105
use FILL  FILL_1376
timestamp 1681708930
transform 1 0 224 0 -1 370
box -8 -3 16 105
use FILL  FILL_1377
timestamp 1681708930
transform 1 0 232 0 -1 370
box -8 -3 16 105
use FILL  FILL_1378
timestamp 1681708930
transform 1 0 240 0 -1 370
box -8 -3 16 105
use FILL  FILL_1379
timestamp 1681708930
transform 1 0 248 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_233
timestamp 1681708930
transform 1 0 256 0 -1 370
box -9 -3 26 105
use OAI21X1  OAI21X1_95
timestamp 1681708930
transform 1 0 272 0 -1 370
box -8 -3 34 105
use FILL  FILL_1380
timestamp 1681708930
transform 1 0 304 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_234
timestamp 1681708930
transform 1 0 312 0 -1 370
box -9 -3 26 105
use FILL  FILL_1381
timestamp 1681708930
transform 1 0 328 0 -1 370
box -8 -3 16 105
use FILL  FILL_1382
timestamp 1681708930
transform 1 0 336 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_235
timestamp 1681708930
transform -1 0 360 0 -1 370
box -9 -3 26 105
use FILL  FILL_1383
timestamp 1681708930
transform 1 0 360 0 -1 370
box -8 -3 16 105
use FILL  FILL_1384
timestamp 1681708930
transform 1 0 368 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_236
timestamp 1681708930
transform -1 0 392 0 -1 370
box -9 -3 26 105
use FILL  FILL_1385
timestamp 1681708930
transform 1 0 392 0 -1 370
box -8 -3 16 105
use FILL  FILL_1386
timestamp 1681708930
transform 1 0 400 0 -1 370
box -8 -3 16 105
use FILL  FILL_1387
timestamp 1681708930
transform 1 0 408 0 -1 370
box -8 -3 16 105
use FILL  FILL_1388
timestamp 1681708930
transform 1 0 416 0 -1 370
box -8 -3 16 105
use FILL  FILL_1389
timestamp 1681708930
transform 1 0 424 0 -1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_96
timestamp 1681708930
transform 1 0 432 0 -1 370
box -8 -3 34 105
use FILL  FILL_1390
timestamp 1681708930
transform 1 0 464 0 -1 370
box -8 -3 16 105
use FILL  FILL_1391
timestamp 1681708930
transform 1 0 472 0 -1 370
box -8 -3 16 105
use FILL  FILL_1392
timestamp 1681708930
transform 1 0 480 0 -1 370
box -8 -3 16 105
use FILL  FILL_1393
timestamp 1681708930
transform 1 0 488 0 -1 370
box -8 -3 16 105
use FILL  FILL_1394
timestamp 1681708930
transform 1 0 496 0 -1 370
box -8 -3 16 105
use FILL  FILL_1395
timestamp 1681708930
transform 1 0 504 0 -1 370
box -8 -3 16 105
use FILL  FILL_1396
timestamp 1681708930
transform 1 0 512 0 -1 370
box -8 -3 16 105
use FILL  FILL_1397
timestamp 1681708930
transform 1 0 520 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_91
timestamp 1681708930
transform 1 0 528 0 -1 370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_92
timestamp 1681708930
transform 1 0 568 0 -1 370
box -8 -3 104 105
use NAND2X1  NAND2X1_84
timestamp 1681708930
transform 1 0 664 0 -1 370
box -8 -3 32 105
use OAI21X1  OAI21X1_97
timestamp 1681708930
transform -1 0 720 0 -1 370
box -8 -3 34 105
use FILL  FILL_1398
timestamp 1681708930
transform 1 0 720 0 -1 370
box -8 -3 16 105
use FILL  FILL_1399
timestamp 1681708930
transform 1 0 728 0 -1 370
box -8 -3 16 105
use FILL  FILL_1400
timestamp 1681708930
transform 1 0 736 0 -1 370
box -8 -3 16 105
use FILL  FILL_1401
timestamp 1681708930
transform 1 0 744 0 -1 370
box -8 -3 16 105
use FILL  FILL_1402
timestamp 1681708930
transform 1 0 752 0 -1 370
box -8 -3 16 105
use FILL  FILL_1403
timestamp 1681708930
transform 1 0 760 0 -1 370
box -8 -3 16 105
use FILL  FILL_1404
timestamp 1681708930
transform 1 0 768 0 -1 370
box -8 -3 16 105
use FILL  FILL_1405
timestamp 1681708930
transform 1 0 776 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_93
timestamp 1681708930
transform 1 0 784 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_237
timestamp 1681708930
transform 1 0 880 0 -1 370
box -9 -3 26 105
use XOR2X1  XOR2X1_186
timestamp 1681708930
transform -1 0 952 0 -1 370
box -8 -3 64 105
use FILL  FILL_1406
timestamp 1681708930
transform 1 0 952 0 -1 370
box -8 -3 16 105
use FILL  FILL_1408
timestamp 1681708930
transform 1 0 960 0 -1 370
box -8 -3 16 105
use FILL  FILL_1420
timestamp 1681708930
transform 1 0 968 0 -1 370
box -8 -3 16 105
use FILL  FILL_1421
timestamp 1681708930
transform 1 0 976 0 -1 370
box -8 -3 16 105
use FILL  FILL_1422
timestamp 1681708930
transform 1 0 984 0 -1 370
box -8 -3 16 105
use FILL  FILL_1423
timestamp 1681708930
transform 1 0 992 0 -1 370
box -8 -3 16 105
use FILL  FILL_1424
timestamp 1681708930
transform 1 0 1000 0 -1 370
box -8 -3 16 105
use FILL  FILL_1425
timestamp 1681708930
transform 1 0 1008 0 -1 370
box -8 -3 16 105
use FILL  FILL_1426
timestamp 1681708930
transform 1 0 1016 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_95
timestamp 1681708930
transform 1 0 1024 0 -1 370
box -8 -3 46 105
use XOR2X1  XOR2X1_188
timestamp 1681708930
transform -1 0 1120 0 -1 370
box -8 -3 64 105
use FILL  FILL_1427
timestamp 1681708930
transform 1 0 1120 0 -1 370
box -8 -3 16 105
use FILL  FILL_1428
timestamp 1681708930
transform 1 0 1128 0 -1 370
box -8 -3 16 105
use XOR2X1  XOR2X1_189
timestamp 1681708930
transform -1 0 1192 0 -1 370
box -8 -3 64 105
use FILL  FILL_1429
timestamp 1681708930
transform 1 0 1192 0 -1 370
box -8 -3 16 105
use FILL  FILL_1430
timestamp 1681708930
transform 1 0 1200 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_3703
timestamp 1681708930
transform 1 0 1244 0 1 275
box -3 -3 3 3
use XOR2X1  XOR2X1_190
timestamp 1681708930
transform 1 0 1208 0 -1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_191
timestamp 1681708930
transform 1 0 1264 0 -1 370
box -8 -3 64 105
use FILL  FILL_1431
timestamp 1681708930
transform 1 0 1320 0 -1 370
box -8 -3 16 105
use FILL  FILL_1454
timestamp 1681708930
transform 1 0 1328 0 -1 370
box -8 -3 16 105
use FILL  FILL_1455
timestamp 1681708930
transform 1 0 1336 0 -1 370
box -8 -3 16 105
use FILL  FILL_1456
timestamp 1681708930
transform 1 0 1344 0 -1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_136
timestamp 1681708930
transform -1 0 1384 0 -1 370
box -8 -3 40 105
use FILL  FILL_1457
timestamp 1681708930
transform 1 0 1384 0 -1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_137
timestamp 1681708930
transform -1 0 1424 0 -1 370
box -8 -3 40 105
use FILL  FILL_1458
timestamp 1681708930
transform 1 0 1424 0 -1 370
box -8 -3 16 105
use FILL  FILL_1459
timestamp 1681708930
transform 1 0 1432 0 -1 370
box -8 -3 16 105
use FILL  FILL_1460
timestamp 1681708930
transform 1 0 1440 0 -1 370
box -8 -3 16 105
use FILL  FILL_1461
timestamp 1681708930
transform 1 0 1448 0 -1 370
box -8 -3 16 105
use FILL  FILL_1462
timestamp 1681708930
transform 1 0 1456 0 -1 370
box -8 -3 16 105
use FILL  FILL_1463
timestamp 1681708930
transform 1 0 1464 0 -1 370
box -8 -3 16 105
use AOI21X1  AOI21X1_50
timestamp 1681708930
transform -1 0 1504 0 -1 370
box -7 -3 39 105
use FILL  FILL_1464
timestamp 1681708930
transform 1 0 1504 0 -1 370
box -8 -3 16 105
use FILL  FILL_1465
timestamp 1681708930
transform 1 0 1512 0 -1 370
box -8 -3 16 105
use FILL  FILL_1466
timestamp 1681708930
transform 1 0 1520 0 -1 370
box -8 -3 16 105
use FILL  FILL_1467
timestamp 1681708930
transform 1 0 1528 0 -1 370
box -8 -3 16 105
use FILL  FILL_1468
timestamp 1681708930
transform 1 0 1536 0 -1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_86
timestamp 1681708930
transform 1 0 1544 0 -1 370
box -8 -3 32 105
use OAI21X1  OAI21X1_100
timestamp 1681708930
transform 1 0 1568 0 -1 370
box -8 -3 34 105
use FILL  FILL_1469
timestamp 1681708930
transform 1 0 1600 0 -1 370
box -8 -3 16 105
use FILL  FILL_1470
timestamp 1681708930
transform 1 0 1608 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_240
timestamp 1681708930
transform 1 0 1616 0 -1 370
box -9 -3 26 105
use NAND2X1  NAND2X1_87
timestamp 1681708930
transform -1 0 1656 0 -1 370
box -8 -3 32 105
use AOI21X1  AOI21X1_51
timestamp 1681708930
transform -1 0 1688 0 -1 370
box -7 -3 39 105
use OAI21X1  OAI21X1_101
timestamp 1681708930
transform -1 0 1720 0 -1 370
box -8 -3 34 105
use XNOR2X1  XNOR2X1_53
timestamp 1681708930
transform 1 0 1720 0 -1 370
box -8 -3 64 105
use FILL  FILL_1471
timestamp 1681708930
transform 1 0 1776 0 -1 370
box -8 -3 16 105
use OR2X1  OR2X1_24
timestamp 1681708930
transform -1 0 1816 0 -1 370
box -8 -3 40 105
use FILL  FILL_1472
timestamp 1681708930
transform 1 0 1816 0 -1 370
box -8 -3 16 105
use FILL  FILL_1473
timestamp 1681708930
transform 1 0 1824 0 -1 370
box -8 -3 16 105
use FILL  FILL_1474
timestamp 1681708930
transform 1 0 1832 0 -1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_138
timestamp 1681708930
transform -1 0 1872 0 -1 370
box -8 -3 40 105
use FILL  FILL_1475
timestamp 1681708930
transform 1 0 1872 0 -1 370
box -8 -3 16 105
use FILL  FILL_1476
timestamp 1681708930
transform 1 0 1880 0 -1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_102
timestamp 1681708930
transform -1 0 1920 0 -1 370
box -8 -3 34 105
use AOI21X1  AOI21X1_52
timestamp 1681708930
transform 1 0 1920 0 -1 370
box -7 -3 39 105
use NOR2X1  NOR2X1_82
timestamp 1681708930
transform -1 0 1976 0 -1 370
box -8 -3 32 105
use INVX2  INVX2_241
timestamp 1681708930
transform -1 0 1992 0 -1 370
box -9 -3 26 105
use NAND3X1  NAND3X1_139
timestamp 1681708930
transform -1 0 2024 0 -1 370
box -8 -3 40 105
use NOR2X1  NOR2X1_83
timestamp 1681708930
transform 1 0 2024 0 -1 370
box -8 -3 32 105
use OAI21X1  OAI21X1_103
timestamp 1681708930
transform -1 0 2080 0 -1 370
box -8 -3 34 105
use INVX2  INVX2_242
timestamp 1681708930
transform 1 0 2080 0 -1 370
box -9 -3 26 105
use M3_M2  M3_M2_3704
timestamp 1681708930
transform 1 0 2140 0 1 275
box -3 -3 3 3
use AOI22X1  AOI22X1_96
timestamp 1681708930
transform 1 0 2096 0 -1 370
box -8 -3 46 105
use FILL  FILL_1477
timestamp 1681708930
transform 1 0 2136 0 -1 370
box -8 -3 16 105
use FILL  FILL_1478
timestamp 1681708930
transform 1 0 2144 0 -1 370
box -8 -3 16 105
use FILL  FILL_1479
timestamp 1681708930
transform 1 0 2152 0 -1 370
box -8 -3 16 105
use FILL  FILL_1480
timestamp 1681708930
transform 1 0 2160 0 -1 370
box -8 -3 16 105
use FILL  FILL_1481
timestamp 1681708930
transform 1 0 2168 0 -1 370
box -8 -3 16 105
use FILL  FILL_1482
timestamp 1681708930
transform 1 0 2176 0 -1 370
box -8 -3 16 105
use OR2X1  OR2X1_25
timestamp 1681708930
transform -1 0 2216 0 -1 370
box -8 -3 40 105
use OAI21X1  OAI21X1_104
timestamp 1681708930
transform -1 0 2248 0 -1 370
box -8 -3 34 105
use INVX2  INVX2_243
timestamp 1681708930
transform 1 0 2248 0 -1 370
box -9 -3 26 105
use NAND3X1  NAND3X1_140
timestamp 1681708930
transform -1 0 2296 0 -1 370
box -8 -3 40 105
use AOI22X1  AOI22X1_97
timestamp 1681708930
transform 1 0 2296 0 -1 370
box -8 -3 46 105
use FILL  FILL_1483
timestamp 1681708930
transform 1 0 2336 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_245
timestamp 1681708930
transform 1 0 2344 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_246
timestamp 1681708930
transform -1 0 2376 0 -1 370
box -9 -3 26 105
use NOR2X1  NOR2X1_85
timestamp 1681708930
transform 1 0 2376 0 -1 370
box -8 -3 32 105
use NAND3X1  NAND3X1_144
timestamp 1681708930
transform 1 0 2400 0 -1 370
box -8 -3 40 105
use INVX2  INVX2_247
timestamp 1681708930
transform -1 0 2448 0 -1 370
box -9 -3 26 105
use FILL  FILL_1489
timestamp 1681708930
transform 1 0 2448 0 -1 370
box -8 -3 16 105
use FILL  FILL_1490
timestamp 1681708930
transform 1 0 2456 0 -1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_90
timestamp 1681708930
transform 1 0 2464 0 -1 370
box -8 -3 32 105
use OAI21X1  OAI21X1_107
timestamp 1681708930
transform -1 0 2520 0 -1 370
box -8 -3 34 105
use NAND2X1  NAND2X1_91
timestamp 1681708930
transform 1 0 2520 0 -1 370
box -8 -3 32 105
use OAI21X1  OAI21X1_108
timestamp 1681708930
transform 1 0 2544 0 -1 370
box -8 -3 34 105
use AOI21X1  AOI21X1_53
timestamp 1681708930
transform -1 0 2608 0 -1 370
box -7 -3 39 105
use XNOR2X1  XNOR2X1_54
timestamp 1681708930
transform -1 0 2664 0 -1 370
box -8 -3 64 105
use top_mod_new_VIA0  top_mod_new_VIA0_47
timestamp 1681708930
transform 1 0 2712 0 1 270
box -10 -3 10 3
use M2_M1  M2_M1_3889
timestamp 1681708930
transform 1 0 76 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3890
timestamp 1681708930
transform 1 0 132 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3861
timestamp 1681708930
transform 1 0 188 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3956
timestamp 1681708930
transform 1 0 156 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3957
timestamp 1681708930
transform 1 0 172 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3958
timestamp 1681708930
transform 1 0 188 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3793
timestamp 1681708930
transform 1 0 68 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3794
timestamp 1681708930
transform 1 0 132 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3795
timestamp 1681708930
transform 1 0 188 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_3891
timestamp 1681708930
transform 1 0 220 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3892
timestamp 1681708930
transform 1 0 228 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3893
timestamp 1681708930
transform 1 0 284 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3959
timestamp 1681708930
transform 1 0 220 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3960
timestamp 1681708930
transform 1 0 308 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3796
timestamp 1681708930
transform 1 0 308 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3705
timestamp 1681708930
transform 1 0 444 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_3723
timestamp 1681708930
transform 1 0 428 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_3862
timestamp 1681708930
transform 1 0 444 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3894
timestamp 1681708930
transform 1 0 380 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3895
timestamp 1681708930
transform 1 0 412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3896
timestamp 1681708930
transform 1 0 428 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3961
timestamp 1681708930
transform 1 0 332 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3962
timestamp 1681708930
transform 1 0 420 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3797
timestamp 1681708930
transform 1 0 332 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3798
timestamp 1681708930
transform 1 0 380 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3706
timestamp 1681708930
transform 1 0 548 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_3707
timestamp 1681708930
transform 1 0 564 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_3897
timestamp 1681708930
transform 1 0 452 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3898
timestamp 1681708930
transform 1 0 508 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3863
timestamp 1681708930
transform 1 0 564 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3963
timestamp 1681708930
transform 1 0 444 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3964
timestamp 1681708930
transform 1 0 532 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3965
timestamp 1681708930
transform 1 0 548 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3966
timestamp 1681708930
transform 1 0 564 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3799
timestamp 1681708930
transform 1 0 444 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3800
timestamp 1681708930
transform 1 0 508 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3801
timestamp 1681708930
transform 1 0 564 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3826
timestamp 1681708930
transform 1 0 452 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3827
timestamp 1681708930
transform 1 0 548 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_3864
timestamp 1681708930
transform 1 0 700 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3899
timestamp 1681708930
transform 1 0 596 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3900
timestamp 1681708930
transform 1 0 660 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3901
timestamp 1681708930
transform 1 0 692 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3967
timestamp 1681708930
transform 1 0 596 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3968
timestamp 1681708930
transform 1 0 612 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3802
timestamp 1681708930
transform 1 0 660 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_3969
timestamp 1681708930
transform 1 0 716 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3970
timestamp 1681708930
transform 1 0 724 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3803
timestamp 1681708930
transform 1 0 724 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3828
timestamp 1681708930
transform 1 0 660 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3829
timestamp 1681708930
transform 1 0 692 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3830
timestamp 1681708930
transform 1 0 716 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3742
timestamp 1681708930
transform 1 0 748 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3724
timestamp 1681708930
transform 1 0 844 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3725
timestamp 1681708930
transform 1 0 876 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_3902
timestamp 1681708930
transform 1 0 748 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3903
timestamp 1681708930
transform 1 0 812 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3971
timestamp 1681708930
transform 1 0 748 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3972
timestamp 1681708930
transform 1 0 764 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3804
timestamp 1681708930
transform 1 0 812 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3743
timestamp 1681708930
transform 1 0 860 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_3904
timestamp 1681708930
transform 1 0 860 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3905
timestamp 1681708930
transform 1 0 876 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3906
timestamp 1681708930
transform 1 0 892 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3865
timestamp 1681708930
transform 1 0 900 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3973
timestamp 1681708930
transform 1 0 892 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3781
timestamp 1681708930
transform 1 0 900 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_3974
timestamp 1681708930
transform 1 0 908 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3805
timestamp 1681708930
transform 1 0 892 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_3975
timestamp 1681708930
transform 1 0 932 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3726
timestamp 1681708930
transform 1 0 964 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_3866
timestamp 1681708930
transform 1 0 964 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3907
timestamp 1681708930
transform 1 0 956 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3760
timestamp 1681708930
transform 1 0 980 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_3908
timestamp 1681708930
transform 1 0 988 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3761
timestamp 1681708930
transform 1 0 1004 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_3909
timestamp 1681708930
transform 1 0 1012 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3976
timestamp 1681708930
transform 1 0 980 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3977
timestamp 1681708930
transform 1 0 996 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3978
timestamp 1681708930
transform 1 0 1004 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3831
timestamp 1681708930
transform 1 0 996 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_3910
timestamp 1681708930
transform 1 0 1020 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3806
timestamp 1681708930
transform 1 0 1012 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3708
timestamp 1681708930
transform 1 0 1068 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_3711
timestamp 1681708930
transform 1 0 1060 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_3727
timestamp 1681708930
transform 1 0 1044 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3744
timestamp 1681708930
transform 1 0 1068 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_3911
timestamp 1681708930
transform 1 0 1044 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3912
timestamp 1681708930
transform 1 0 1060 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3782
timestamp 1681708930
transform 1 0 1044 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_3979
timestamp 1681708930
transform 1 0 1052 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3832
timestamp 1681708930
transform 1 0 1052 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_3980
timestamp 1681708930
transform 1 0 1068 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3913
timestamp 1681708930
transform 1 0 1084 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3745
timestamp 1681708930
transform 1 0 1220 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_3914
timestamp 1681708930
transform 1 0 1164 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3981
timestamp 1681708930
transform 1 0 1132 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3982
timestamp 1681708930
transform 1 0 1140 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3807
timestamp 1681708930
transform 1 0 1140 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3762
timestamp 1681708930
transform 1 0 1196 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_3915
timestamp 1681708930
transform 1 0 1220 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3983
timestamp 1681708930
transform 1 0 1196 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3984
timestamp 1681708930
transform 1 0 1244 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3985
timestamp 1681708930
transform 1 0 1252 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3712
timestamp 1681708930
transform 1 0 1292 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_3916
timestamp 1681708930
transform 1 0 1292 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3808
timestamp 1681708930
transform 1 0 1268 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3709
timestamp 1681708930
transform 1 0 1332 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_3867
timestamp 1681708930
transform 1 0 1324 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_3763
timestamp 1681708930
transform 1 0 1324 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_3986
timestamp 1681708930
transform 1 0 1332 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3746
timestamp 1681708930
transform 1 0 1356 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_3917
timestamp 1681708930
transform 1 0 1356 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3717
timestamp 1681708930
transform 1 0 1380 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_3854
timestamp 1681708930
transform 1 0 1380 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_4024
timestamp 1681708930
transform 1 0 1380 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_3747
timestamp 1681708930
transform 1 0 1412 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_3868
timestamp 1681708930
transform 1 0 1420 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_3713
timestamp 1681708930
transform 1 0 1444 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_3855
timestamp 1681708930
transform 1 0 1452 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_3869
timestamp 1681708930
transform 1 0 1444 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3870
timestamp 1681708930
transform 1 0 1452 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3918
timestamp 1681708930
transform 1 0 1412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3919
timestamp 1681708930
transform 1 0 1436 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3987
timestamp 1681708930
transform 1 0 1404 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3809
timestamp 1681708930
transform 1 0 1404 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3764
timestamp 1681708930
transform 1 0 1452 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_3714
timestamp 1681708930
transform 1 0 1508 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_3728
timestamp 1681708930
transform 1 0 1484 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_3856
timestamp 1681708930
transform 1 0 1500 0 1 235
box -2 -2 2 2
use M3_M2  M3_M2_3748
timestamp 1681708930
transform 1 0 1476 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_3871
timestamp 1681708930
transform 1 0 1492 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3988
timestamp 1681708930
transform 1 0 1460 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3920
timestamp 1681708930
transform 1 0 1484 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3765
timestamp 1681708930
transform 1 0 1492 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_3921
timestamp 1681708930
transform 1 0 1508 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3989
timestamp 1681708930
transform 1 0 1484 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3783
timestamp 1681708930
transform 1 0 1500 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_3872
timestamp 1681708930
transform 1 0 1524 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_3749
timestamp 1681708930
transform 1 0 1532 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_3922
timestamp 1681708930
transform 1 0 1524 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3766
timestamp 1681708930
transform 1 0 1532 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_3990
timestamp 1681708930
transform 1 0 1532 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3810
timestamp 1681708930
transform 1 0 1524 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3715
timestamp 1681708930
transform 1 0 1588 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_3729
timestamp 1681708930
transform 1 0 1572 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3716
timestamp 1681708930
transform 1 0 1628 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_3730
timestamp 1681708930
transform 1 0 1628 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3750
timestamp 1681708930
transform 1 0 1564 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3751
timestamp 1681708930
transform 1 0 1596 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3752
timestamp 1681708930
transform 1 0 1620 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_3923
timestamp 1681708930
transform 1 0 1572 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3924
timestamp 1681708930
transform 1 0 1588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3925
timestamp 1681708930
transform 1 0 1596 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3991
timestamp 1681708930
transform 1 0 1564 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3992
timestamp 1681708930
transform 1 0 1588 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3993
timestamp 1681708930
transform 1 0 1596 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3811
timestamp 1681708930
transform 1 0 1588 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3784
timestamp 1681708930
transform 1 0 1604 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_3926
timestamp 1681708930
transform 1 0 1628 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3994
timestamp 1681708930
transform 1 0 1620 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3995
timestamp 1681708930
transform 1 0 1628 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3833
timestamp 1681708930
transform 1 0 1604 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3731
timestamp 1681708930
transform 1 0 1652 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_3857
timestamp 1681708930
transform 1 0 1668 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_3873
timestamp 1681708930
transform 1 0 1652 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3874
timestamp 1681708930
transform 1 0 1660 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_3753
timestamp 1681708930
transform 1 0 1668 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_3875
timestamp 1681708930
transform 1 0 1684 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3927
timestamp 1681708930
transform 1 0 1652 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3928
timestamp 1681708930
transform 1 0 1676 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3812
timestamp 1681708930
transform 1 0 1644 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3834
timestamp 1681708930
transform 1 0 1628 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3767
timestamp 1681708930
transform 1 0 1684 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_3813
timestamp 1681708930
transform 1 0 1676 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3768
timestamp 1681708930
transform 1 0 1700 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_3996
timestamp 1681708930
transform 1 0 1700 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3718
timestamp 1681708930
transform 1 0 1716 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_3929
timestamp 1681708930
transform 1 0 1708 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3930
timestamp 1681708930
transform 1 0 1716 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3769
timestamp 1681708930
transform 1 0 1732 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_3997
timestamp 1681708930
transform 1 0 1732 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4025
timestamp 1681708930
transform 1 0 1716 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_3835
timestamp 1681708930
transform 1 0 1724 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3732
timestamp 1681708930
transform 1 0 1748 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_3931
timestamp 1681708930
transform 1 0 1748 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3836
timestamp 1681708930
transform 1 0 1748 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3710
timestamp 1681708930
transform 1 0 1772 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_3785
timestamp 1681708930
transform 1 0 1780 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_3814
timestamp 1681708930
transform 1 0 1772 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_4026
timestamp 1681708930
transform 1 0 1780 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_3998
timestamp 1681708930
transform 1 0 1820 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3770
timestamp 1681708930
transform 1 0 1844 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_3932
timestamp 1681708930
transform 1 0 1852 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3999
timestamp 1681708930
transform 1 0 1836 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4027
timestamp 1681708930
transform 1 0 1828 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_3786
timestamp 1681708930
transform 1 0 1852 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_4028
timestamp 1681708930
transform 1 0 1852 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_3933
timestamp 1681708930
transform 1 0 1868 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3733
timestamp 1681708930
transform 1 0 1892 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_3934
timestamp 1681708930
transform 1 0 1892 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3771
timestamp 1681708930
transform 1 0 1900 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_4000
timestamp 1681708930
transform 1 0 1940 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3719
timestamp 1681708930
transform 1 0 1956 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_3734
timestamp 1681708930
transform 1 0 1996 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_3876
timestamp 1681708930
transform 1 0 1956 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_3754
timestamp 1681708930
transform 1 0 1972 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3772
timestamp 1681708930
transform 1 0 1956 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_3935
timestamp 1681708930
transform 1 0 1972 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3773
timestamp 1681708930
transform 1 0 1980 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_3936
timestamp 1681708930
transform 1 0 1988 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3787
timestamp 1681708930
transform 1 0 1980 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_4001
timestamp 1681708930
transform 1 0 1988 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3877
timestamp 1681708930
transform 1 0 1996 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_3755
timestamp 1681708930
transform 1 0 2020 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_3878
timestamp 1681708930
transform 1 0 2028 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3937
timestamp 1681708930
transform 1 0 2012 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3938
timestamp 1681708930
transform 1 0 2020 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3774
timestamp 1681708930
transform 1 0 2028 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_4002
timestamp 1681708930
transform 1 0 2028 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3735
timestamp 1681708930
transform 1 0 2044 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_3879
timestamp 1681708930
transform 1 0 2044 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_3720
timestamp 1681708930
transform 1 0 2060 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_3858
timestamp 1681708930
transform 1 0 2068 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_3880
timestamp 1681708930
transform 1 0 2076 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4003
timestamp 1681708930
transform 1 0 2052 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3788
timestamp 1681708930
transform 1 0 2060 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_4004
timestamp 1681708930
transform 1 0 2076 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3789
timestamp 1681708930
transform 1 0 2084 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_4005
timestamp 1681708930
transform 1 0 2092 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3815
timestamp 1681708930
transform 1 0 2076 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3837
timestamp 1681708930
transform 1 0 2092 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3721
timestamp 1681708930
transform 1 0 2108 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_3939
timestamp 1681708930
transform 1 0 2100 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3940
timestamp 1681708930
transform 1 0 2108 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4006
timestamp 1681708930
transform 1 0 2108 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3816
timestamp 1681708930
transform 1 0 2108 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3756
timestamp 1681708930
transform 1 0 2124 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_3941
timestamp 1681708930
transform 1 0 2124 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4007
timestamp 1681708930
transform 1 0 2124 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3838
timestamp 1681708930
transform 1 0 2124 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3722
timestamp 1681708930
transform 1 0 2172 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_3736
timestamp 1681708930
transform 1 0 2196 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_3859
timestamp 1681708930
transform 1 0 2204 0 1 235
box -2 -2 2 2
use M3_M2  M3_M2_3737
timestamp 1681708930
transform 1 0 2228 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_3860
timestamp 1681708930
transform 1 0 2244 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_3881
timestamp 1681708930
transform 1 0 2180 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3882
timestamp 1681708930
transform 1 0 2204 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3883
timestamp 1681708930
transform 1 0 2228 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3942
timestamp 1681708930
transform 1 0 2196 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4008
timestamp 1681708930
transform 1 0 2172 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3775
timestamp 1681708930
transform 1 0 2204 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_3943
timestamp 1681708930
transform 1 0 2212 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3790
timestamp 1681708930
transform 1 0 2212 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_3738
timestamp 1681708930
transform 1 0 2252 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3739
timestamp 1681708930
transform 1 0 2276 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_3884
timestamp 1681708930
transform 1 0 2252 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3944
timestamp 1681708930
transform 1 0 2244 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4009
timestamp 1681708930
transform 1 0 2220 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3817
timestamp 1681708930
transform 1 0 2228 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3839
timestamp 1681708930
transform 1 0 2220 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_3885
timestamp 1681708930
transform 1 0 2284 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_3776
timestamp 1681708930
transform 1 0 2284 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_4010
timestamp 1681708930
transform 1 0 2268 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4011
timestamp 1681708930
transform 1 0 2276 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4012
timestamp 1681708930
transform 1 0 2284 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4029
timestamp 1681708930
transform 1 0 2260 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_3945
timestamp 1681708930
transform 1 0 2316 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3777
timestamp 1681708930
transform 1 0 2324 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_3946
timestamp 1681708930
transform 1 0 2332 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3947
timestamp 1681708930
transform 1 0 2340 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4013
timestamp 1681708930
transform 1 0 2308 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3791
timestamp 1681708930
transform 1 0 2340 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_3740
timestamp 1681708930
transform 1 0 2412 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3741
timestamp 1681708930
transform 1 0 2428 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3757
timestamp 1681708930
transform 1 0 2372 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3758
timestamp 1681708930
transform 1 0 2404 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3778
timestamp 1681708930
transform 1 0 2364 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_3948
timestamp 1681708930
transform 1 0 2372 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3949
timestamp 1681708930
transform 1 0 2404 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4014
timestamp 1681708930
transform 1 0 2356 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4015
timestamp 1681708930
transform 1 0 2364 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3818
timestamp 1681708930
transform 1 0 2308 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_4030
timestamp 1681708930
transform 1 0 2316 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_3819
timestamp 1681708930
transform 1 0 2324 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_4031
timestamp 1681708930
transform 1 0 2332 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_3820
timestamp 1681708930
transform 1 0 2356 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3840
timestamp 1681708930
transform 1 0 2332 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_4016
timestamp 1681708930
transform 1 0 2420 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4017
timestamp 1681708930
transform 1 0 2428 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3821
timestamp 1681708930
transform 1 0 2428 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3759
timestamp 1681708930
transform 1 0 2436 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_3950
timestamp 1681708930
transform 1 0 2436 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3951
timestamp 1681708930
transform 1 0 2444 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4018
timestamp 1681708930
transform 1 0 2460 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4032
timestamp 1681708930
transform 1 0 2444 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_3822
timestamp 1681708930
transform 1 0 2460 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_3886
timestamp 1681708930
transform 1 0 2516 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3887
timestamp 1681708930
transform 1 0 2540 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3888
timestamp 1681708930
transform 1 0 2548 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3952
timestamp 1681708930
transform 1 0 2492 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3953
timestamp 1681708930
transform 1 0 2508 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_3792
timestamp 1681708930
transform 1 0 2484 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_4019
timestamp 1681708930
transform 1 0 2492 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4033
timestamp 1681708930
transform 1 0 2476 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_3841
timestamp 1681708930
transform 1 0 2444 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3823
timestamp 1681708930
transform 1 0 2484 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3779
timestamp 1681708930
transform 1 0 2516 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_3780
timestamp 1681708930
transform 1 0 2540 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_3954
timestamp 1681708930
transform 1 0 2548 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3955
timestamp 1681708930
transform 1 0 2564 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4020
timestamp 1681708930
transform 1 0 2516 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4021
timestamp 1681708930
transform 1 0 2540 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3842
timestamp 1681708930
transform 1 0 2540 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_4022
timestamp 1681708930
transform 1 0 2580 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3824
timestamp 1681708930
transform 1 0 2580 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_4023
timestamp 1681708930
transform 1 0 2628 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_3825
timestamp 1681708930
transform 1 0 2628 0 1 195
box -3 -3 3 3
use top_mod_new_VIA0  top_mod_new_VIA0_48
timestamp 1681708930
transform 1 0 48 0 1 170
box -10 -3 10 3
use M3_M2  M3_M2_3843
timestamp 1681708930
transform 1 0 76 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3844
timestamp 1681708930
transform 1 0 172 0 1 175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_94
timestamp 1681708930
transform -1 0 168 0 1 170
box -8 -3 104 105
use NAND2X1  NAND2X1_92
timestamp 1681708930
transform 1 0 168 0 1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_109
timestamp 1681708930
transform -1 0 224 0 1 170
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_95
timestamp 1681708930
transform -1 0 320 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_96
timestamp 1681708930
transform 1 0 320 0 1 170
box -8 -3 104 105
use OAI21X1  OAI21X1_110
timestamp 1681708930
transform 1 0 416 0 1 170
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_97
timestamp 1681708930
transform -1 0 544 0 1 170
box -8 -3 104 105
use NAND2X1  NAND2X1_93
timestamp 1681708930
transform 1 0 544 0 1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_111
timestamp 1681708930
transform -1 0 600 0 1 170
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_98
timestamp 1681708930
transform 1 0 600 0 1 170
box -8 -3 104 105
use NAND2X1  NAND2X1_94
timestamp 1681708930
transform -1 0 720 0 1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_112
timestamp 1681708930
transform -1 0 752 0 1 170
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_99
timestamp 1681708930
transform 1 0 752 0 1 170
box -8 -3 104 105
use INVX2  INVX2_248
timestamp 1681708930
transform 1 0 848 0 1 170
box -9 -3 26 105
use OAI21X1  OAI21X1_113
timestamp 1681708930
transform 1 0 864 0 1 170
box -8 -3 34 105
use FILL  FILL_1491
timestamp 1681708930
transform 1 0 896 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_114
timestamp 1681708930
transform 1 0 904 0 1 170
box -8 -3 34 105
use FILL  FILL_1492
timestamp 1681708930
transform 1 0 936 0 1 170
box -8 -3 16 105
use FILL  FILL_1493
timestamp 1681708930
transform 1 0 944 0 1 170
box -8 -3 16 105
use FILL  FILL_1494
timestamp 1681708930
transform 1 0 952 0 1 170
box -8 -3 16 105
use FILL  FILL_1495
timestamp 1681708930
transform 1 0 960 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_98
timestamp 1681708930
transform 1 0 968 0 1 170
box -8 -3 46 105
use FILL  FILL_1496
timestamp 1681708930
transform 1 0 1008 0 1 170
box -8 -3 16 105
use FILL  FILL_1497
timestamp 1681708930
transform 1 0 1016 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_99
timestamp 1681708930
transform 1 0 1024 0 1 170
box -8 -3 46 105
use FILL  FILL_1498
timestamp 1681708930
transform 1 0 1064 0 1 170
box -8 -3 16 105
use FILL  FILL_1499
timestamp 1681708930
transform 1 0 1072 0 1 170
box -8 -3 16 105
use XOR2X1  XOR2X1_199
timestamp 1681708930
transform -1 0 1136 0 1 170
box -8 -3 64 105
use XOR2X1  XOR2X1_200
timestamp 1681708930
transform -1 0 1192 0 1 170
box -8 -3 64 105
use XOR2X1  XOR2X1_201
timestamp 1681708930
transform 1 0 1192 0 1 170
box -8 -3 64 105
use FILL  FILL_1500
timestamp 1681708930
transform 1 0 1248 0 1 170
box -8 -3 16 105
use FILL  FILL_1501
timestamp 1681708930
transform 1 0 1256 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_3845
timestamp 1681708930
transform 1 0 1276 0 1 175
box -3 -3 3 3
use XOR2X1  XOR2X1_202
timestamp 1681708930
transform 1 0 1264 0 1 170
box -8 -3 64 105
use FILL  FILL_1502
timestamp 1681708930
transform 1 0 1320 0 1 170
box -8 -3 16 105
use FILL  FILL_1503
timestamp 1681708930
transform 1 0 1328 0 1 170
box -8 -3 16 105
use NAND3X1  NAND3X1_145
timestamp 1681708930
transform -1 0 1368 0 1 170
box -8 -3 40 105
use FILL  FILL_1504
timestamp 1681708930
transform 1 0 1368 0 1 170
box -8 -3 16 105
use FILL  FILL_1505
timestamp 1681708930
transform 1 0 1376 0 1 170
box -8 -3 16 105
use AOI21X1  AOI21X1_54
timestamp 1681708930
transform -1 0 1416 0 1 170
box -7 -3 39 105
use NAND3X1  NAND3X1_146
timestamp 1681708930
transform -1 0 1448 0 1 170
box -8 -3 40 105
use M3_M2  M3_M2_3846
timestamp 1681708930
transform 1 0 1460 0 1 175
box -3 -3 3 3
use FILL  FILL_1506
timestamp 1681708930
transform 1 0 1448 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_115
timestamp 1681708930
transform -1 0 1488 0 1 170
box -8 -3 34 105
use NAND3X1  NAND3X1_147
timestamp 1681708930
transform -1 0 1520 0 1 170
box -8 -3 40 105
use FILL  FILL_1507
timestamp 1681708930
transform 1 0 1520 0 1 170
box -8 -3 16 105
use INVX2  INVX2_253
timestamp 1681708930
transform 1 0 1528 0 1 170
box -9 -3 26 105
use FILL  FILL_1512
timestamp 1681708930
transform 1 0 1544 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_100
timestamp 1681708930
transform 1 0 1552 0 1 170
box -8 -3 46 105
use INVX2  INVX2_254
timestamp 1681708930
transform 1 0 1592 0 1 170
box -9 -3 26 105
use NOR2X1  NOR2X1_88
timestamp 1681708930
transform 1 0 1608 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_99
timestamp 1681708930
transform 1 0 1632 0 1 170
box -8 -3 32 105
use NAND3X1  NAND3X1_150
timestamp 1681708930
transform -1 0 1688 0 1 170
box -8 -3 40 105
use FILL  FILL_1513
timestamp 1681708930
transform 1 0 1688 0 1 170
box -8 -3 16 105
use INVX2  INVX2_255
timestamp 1681708930
transform 1 0 1696 0 1 170
box -9 -3 26 105
use AOI21X1  AOI21X1_56
timestamp 1681708930
transform -1 0 1744 0 1 170
box -7 -3 39 105
use FILL  FILL_1521
timestamp 1681708930
transform 1 0 1744 0 1 170
box -8 -3 16 105
use FILL  FILL_1522
timestamp 1681708930
transform 1 0 1752 0 1 170
box -8 -3 16 105
use NOR2X1  NOR2X1_89
timestamp 1681708930
transform -1 0 1784 0 1 170
box -8 -3 32 105
use FILL  FILL_1523
timestamp 1681708930
transform 1 0 1784 0 1 170
box -8 -3 16 105
use FILL  FILL_1524
timestamp 1681708930
transform 1 0 1792 0 1 170
box -8 -3 16 105
use FILL  FILL_1525
timestamp 1681708930
transform 1 0 1800 0 1 170
box -8 -3 16 105
use FILL  FILL_1526
timestamp 1681708930
transform 1 0 1808 0 1 170
box -8 -3 16 105
use FILL  FILL_1527
timestamp 1681708930
transform 1 0 1816 0 1 170
box -8 -3 16 105
use FILL  FILL_1528
timestamp 1681708930
transform 1 0 1824 0 1 170
box -8 -3 16 105
use INVX2  INVX2_256
timestamp 1681708930
transform 1 0 1832 0 1 170
box -9 -3 26 105
use FILL  FILL_1529
timestamp 1681708930
transform 1 0 1848 0 1 170
box -8 -3 16 105
use FILL  FILL_1534
timestamp 1681708930
transform 1 0 1856 0 1 170
box -8 -3 16 105
use AOI21X1  AOI21X1_57
timestamp 1681708930
transform -1 0 1896 0 1 170
box -7 -3 39 105
use FILL  FILL_1535
timestamp 1681708930
transform 1 0 1896 0 1 170
box -8 -3 16 105
use FILL  FILL_1536
timestamp 1681708930
transform 1 0 1904 0 1 170
box -8 -3 16 105
use FILL  FILL_1537
timestamp 1681708930
transform 1 0 1912 0 1 170
box -8 -3 16 105
use FILL  FILL_1538
timestamp 1681708930
transform 1 0 1920 0 1 170
box -8 -3 16 105
use FILL  FILL_1539
timestamp 1681708930
transform 1 0 1928 0 1 170
box -8 -3 16 105
use NAND2X1  NAND2X1_102
timestamp 1681708930
transform 1 0 1936 0 1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_124
timestamp 1681708930
transform 1 0 1960 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_125
timestamp 1681708930
transform -1 0 2024 0 1 170
box -8 -3 34 105
use NAND2X1  NAND2X1_103
timestamp 1681708930
transform -1 0 2048 0 1 170
box -8 -3 32 105
use FILL  FILL_1540
timestamp 1681708930
transform 1 0 2048 0 1 170
box -8 -3 16 105
use NAND3X1  NAND3X1_151
timestamp 1681708930
transform -1 0 2088 0 1 170
box -8 -3 40 105
use INVX2  INVX2_258
timestamp 1681708930
transform 1 0 2088 0 1 170
box -9 -3 26 105
use INVX2  INVX2_259
timestamp 1681708930
transform 1 0 2104 0 1 170
box -9 -3 26 105
use XNOR2X1  XNOR2X1_57
timestamp 1681708930
transform -1 0 2176 0 1 170
box -8 -3 64 105
use NAND3X1  NAND3X1_152
timestamp 1681708930
transform -1 0 2208 0 1 170
box -8 -3 40 105
use INVX2  INVX2_260
timestamp 1681708930
transform -1 0 2224 0 1 170
box -9 -3 26 105
use NAND3X1  NAND3X1_153
timestamp 1681708930
transform -1 0 2256 0 1 170
box -8 -3 40 105
use M3_M2  M3_M2_3847
timestamp 1681708930
transform 1 0 2284 0 1 175
box -3 -3 3 3
use NOR2X1  NOR2X1_90
timestamp 1681708930
transform 1 0 2256 0 1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_126
timestamp 1681708930
transform -1 0 2312 0 1 170
box -8 -3 34 105
use NOR2X1  NOR2X1_91
timestamp 1681708930
transform 1 0 2312 0 1 170
box -8 -3 32 105
use AOI21X1  AOI21X1_58
timestamp 1681708930
transform -1 0 2368 0 1 170
box -7 -3 39 105
use XNOR2X1  XNOR2X1_58
timestamp 1681708930
transform 1 0 2368 0 1 170
box -8 -3 64 105
use M3_M2  M3_M2_3848
timestamp 1681708930
transform 1 0 2436 0 1 175
box -3 -3 3 3
use INVX2  INVX2_261
timestamp 1681708930
transform 1 0 2424 0 1 170
box -9 -3 26 105
use AOI21X1  AOI21X1_59
timestamp 1681708930
transform -1 0 2472 0 1 170
box -7 -3 39 105
use NOR2X1  NOR2X1_92
timestamp 1681708930
transform 1 0 2472 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_104
timestamp 1681708930
transform 1 0 2496 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_105
timestamp 1681708930
transform 1 0 2520 0 1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_127
timestamp 1681708930
transform -1 0 2576 0 1 170
box -8 -3 34 105
use XNOR2X1  XNOR2X1_59
timestamp 1681708930
transform -1 0 2632 0 1 170
box -8 -3 64 105
use FILL  FILL_1541
timestamp 1681708930
transform 1 0 2632 0 1 170
box -8 -3 16 105
use FILL  FILL_1613
timestamp 1681708930
transform 1 0 2640 0 1 170
box -8 -3 16 105
use FILL  FILL_1615
timestamp 1681708930
transform 1 0 2648 0 1 170
box -8 -3 16 105
use FILL  FILL_1617
timestamp 1681708930
transform 1 0 2656 0 1 170
box -8 -3 16 105
use top_mod_new_VIA0  top_mod_new_VIA0_49
timestamp 1681708930
transform 1 0 2688 0 1 170
box -10 -3 10 3
use M2_M1  M2_M1_4034
timestamp 1681708930
transform 1 0 68 0 1 145
box -2 -2 2 2
use top_mod_new_VIA0  top_mod_new_VIA0_50
timestamp 1681708930
transform 1 0 24 0 1 70
box -10 -3 10 3
use INVX1  INVX1_0
timestamp 1681708930
transform 1 0 72 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_3865
timestamp 1681708930
transform 1 0 156 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3878
timestamp 1681708930
transform 1 0 108 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3879
timestamp 1681708930
transform 1 0 124 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3880
timestamp 1681708930
transform 1 0 156 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3881
timestamp 1681708930
transform 1 0 172 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_4040
timestamp 1681708930
transform 1 0 124 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_3849
timestamp 1681708930
transform 1 0 220 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3882
timestamp 1681708930
transform 1 0 228 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_4041
timestamp 1681708930
transform 1 0 228 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4090
timestamp 1681708930
transform 1 0 108 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4091
timestamp 1681708930
transform 1 0 172 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4092
timestamp 1681708930
transform 1 0 204 0 1 125
box -2 -2 2 2
use INVX4  INVX4_0
timestamp 1681708930
transform 1 0 88 0 -1 170
box -9 -3 28 105
use DFFNEGX1  DFFNEGX1_100
timestamp 1681708930
transform 1 0 112 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_3919
timestamp 1681708930
transform 1 0 228 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3850
timestamp 1681708930
transform 1 0 260 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3866
timestamp 1681708930
transform 1 0 276 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3883
timestamp 1681708930
transform 1 0 324 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_4042
timestamp 1681708930
transform 1 0 260 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4043
timestamp 1681708930
transform 1 0 276 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4093
timestamp 1681708930
transform 1 0 252 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4131
timestamp 1681708930
transform 1 0 228 0 1 115
box -2 -2 2 2
use NAND2X1  NAND2X1_95
timestamp 1681708930
transform 1 0 208 0 -1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_116
timestamp 1681708930
transform -1 0 264 0 -1 170
box -8 -3 34 105
use M3_M2  M3_M2_3884
timestamp 1681708930
transform 1 0 380 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_4044
timestamp 1681708930
transform 1 0 380 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4094
timestamp 1681708930
transform 1 0 324 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4095
timestamp 1681708930
transform 1 0 356 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_3920
timestamp 1681708930
transform 1 0 380 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3851
timestamp 1681708930
transform 1 0 412 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3867
timestamp 1681708930
transform 1 0 428 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3885
timestamp 1681708930
transform 1 0 476 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_4045
timestamp 1681708930
transform 1 0 412 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4046
timestamp 1681708930
transform 1 0 428 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4096
timestamp 1681708930
transform 1 0 404 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4132
timestamp 1681708930
transform 1 0 380 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_3957
timestamp 1681708930
transform 1 0 292 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_3958
timestamp 1681708930
transform 1 0 356 0 1 95
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_101
timestamp 1681708930
transform 1 0 264 0 -1 170
box -8 -3 104 105
use NAND2X1  NAND2X1_96
timestamp 1681708930
transform 1 0 360 0 -1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_117
timestamp 1681708930
transform -1 0 416 0 -1 170
box -8 -3 34 105
use M3_M2  M3_M2_3868
timestamp 1681708930
transform 1 0 532 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3886
timestamp 1681708930
transform 1 0 532 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_4047
timestamp 1681708930
transform 1 0 532 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_3852
timestamp 1681708930
transform 1 0 564 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3853
timestamp 1681708930
transform 1 0 612 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3869
timestamp 1681708930
transform 1 0 580 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3870
timestamp 1681708930
transform 1 0 596 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3887
timestamp 1681708930
transform 1 0 564 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3888
timestamp 1681708930
transform 1 0 596 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3889
timestamp 1681708930
transform 1 0 628 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_4048
timestamp 1681708930
transform 1 0 564 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4049
timestamp 1681708930
transform 1 0 580 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4097
timestamp 1681708930
transform 1 0 476 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4098
timestamp 1681708930
transform 1 0 508 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_3921
timestamp 1681708930
transform 1 0 532 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3922
timestamp 1681708930
transform 1 0 556 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3890
timestamp 1681708930
transform 1 0 684 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_4050
timestamp 1681708930
transform 1 0 684 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_3854
timestamp 1681708930
transform 1 0 764 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3855
timestamp 1681708930
transform 1 0 796 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3871
timestamp 1681708930
transform 1 0 716 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3872
timestamp 1681708930
transform 1 0 748 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3905
timestamp 1681708930
transform 1 0 708 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_3891
timestamp 1681708930
transform 1 0 732 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3892
timestamp 1681708930
transform 1 0 764 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3893
timestamp 1681708930
transform 1 0 780 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_4051
timestamp 1681708930
transform 1 0 716 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4052
timestamp 1681708930
transform 1 0 732 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4099
timestamp 1681708930
transform 1 0 564 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4100
timestamp 1681708930
transform 1 0 628 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4101
timestamp 1681708930
transform 1 0 668 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_3938
timestamp 1681708930
transform 1 0 476 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_3939
timestamp 1681708930
transform 1 0 508 0 1 115
box -3 -3 3 3
use M2_M1  M2_M1_4133
timestamp 1681708930
transform 1 0 532 0 1 115
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_102
timestamp 1681708930
transform 1 0 416 0 -1 170
box -8 -3 104 105
use NAND2X1  NAND2X1_97
timestamp 1681708930
transform 1 0 512 0 -1 170
box -8 -3 32 105
use M3_M2  M3_M2_3940
timestamp 1681708930
transform 1 0 564 0 1 115
box -3 -3 3 3
use OAI21X1  OAI21X1_118
timestamp 1681708930
transform -1 0 568 0 -1 170
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_103
timestamp 1681708930
transform 1 0 568 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_3923
timestamp 1681708930
transform 1 0 684 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3924
timestamp 1681708930
transform 1 0 700 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_4102
timestamp 1681708930
transform 1 0 708 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4134
timestamp 1681708930
transform 1 0 684 0 1 115
box -2 -2 2 2
use NAND2X1  NAND2X1_98
timestamp 1681708930
transform 1 0 664 0 -1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_119
timestamp 1681708930
transform -1 0 720 0 -1 170
box -8 -3 34 105
use M2_M1  M2_M1_4103
timestamp 1681708930
transform 1 0 780 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_104
timestamp 1681708930
transform 1 0 720 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_3873
timestamp 1681708930
transform 1 0 852 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3856
timestamp 1681708930
transform 1 0 876 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3894
timestamp 1681708930
transform 1 0 860 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_4053
timestamp 1681708930
transform 1 0 860 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4054
timestamp 1681708930
transform 1 0 876 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4104
timestamp 1681708930
transform 1 0 828 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4105
timestamp 1681708930
transform 1 0 844 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_3941
timestamp 1681708930
transform 1 0 828 0 1 115
box -3 -3 3 3
use INVX2  INVX2_249
timestamp 1681708930
transform 1 0 816 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_3906
timestamp 1681708930
transform 1 0 908 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_4106
timestamp 1681708930
transform 1 0 924 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4135
timestamp 1681708930
transform 1 0 860 0 1 115
box -2 -2 2 2
use OAI21X1  OAI21X1_120
timestamp 1681708930
transform 1 0 832 0 -1 170
box -8 -3 34 105
use M3_M2  M3_M2_3942
timestamp 1681708930
transform 1 0 948 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_105
timestamp 1681708930
transform 1 0 864 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_3857
timestamp 1681708930
transform 1 0 1028 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3874
timestamp 1681708930
transform 1 0 988 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3907
timestamp 1681708930
transform 1 0 972 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_4055
timestamp 1681708930
transform 1 0 980 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_3875
timestamp 1681708930
transform 1 0 1060 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_4056
timestamp 1681708930
transform 1 0 1028 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4057
timestamp 1681708930
transform 1 0 1036 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4107
timestamp 1681708930
transform 1 0 972 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4108
timestamp 1681708930
transform 1 0 996 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_3943
timestamp 1681708930
transform 1 0 996 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_3947
timestamp 1681708930
transform 1 0 980 0 1 105
box -3 -3 3 3
use INVX2  INVX2_250
timestamp 1681708930
transform 1 0 960 0 -1 170
box -9 -3 26 105
use M2_M1  M2_M1_4058
timestamp 1681708930
transform 1 0 1092 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4109
timestamp 1681708930
transform 1 0 1060 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_3944
timestamp 1681708930
transform 1 0 1060 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_3959
timestamp 1681708930
transform 1 0 1036 0 1 95
box -3 -3 3 3
use XOR2X1  XOR2X1_203
timestamp 1681708930
transform -1 0 1032 0 -1 170
box -8 -3 64 105
use M3_M2  M3_M2_3876
timestamp 1681708930
transform 1 0 1148 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3895
timestamp 1681708930
transform 1 0 1140 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_4059
timestamp 1681708930
transform 1 0 1140 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4060
timestamp 1681708930
transform 1 0 1148 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4110
timestamp 1681708930
transform 1 0 1116 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_3948
timestamp 1681708930
transform 1 0 1116 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_3963
timestamp 1681708930
transform 1 0 1092 0 1 75
box -3 -3 3 3
use XOR2X1  XOR2X1_204
timestamp 1681708930
transform -1 0 1088 0 -1 170
box -8 -3 64 105
use XOR2X1  XOR2X1_205
timestamp 1681708930
transform 1 0 1088 0 -1 170
box -8 -3 64 105
use M3_M2  M3_M2_3858
timestamp 1681708930
transform 1 0 1204 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_4061
timestamp 1681708930
transform 1 0 1196 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4062
timestamp 1681708930
transform 1 0 1204 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4111
timestamp 1681708930
transform 1 0 1172 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_3949
timestamp 1681708930
transform 1 0 1196 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_3960
timestamp 1681708930
transform 1 0 1172 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_3961
timestamp 1681708930
transform 1 0 1204 0 1 95
box -3 -3 3 3
use XOR2X1  XOR2X1_206
timestamp 1681708930
transform 1 0 1144 0 -1 170
box -8 -3 64 105
use M3_M2  M3_M2_3859
timestamp 1681708930
transform 1 0 1252 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3896
timestamp 1681708930
transform 1 0 1260 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3897
timestamp 1681708930
transform 1 0 1292 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_4063
timestamp 1681708930
transform 1 0 1252 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4064
timestamp 1681708930
transform 1 0 1276 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4065
timestamp 1681708930
transform 1 0 1292 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4112
timestamp 1681708930
transform 1 0 1252 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4113
timestamp 1681708930
transform 1 0 1260 0 1 125
box -2 -2 2 2
use XOR2X1  XOR2X1_207
timestamp 1681708930
transform 1 0 1200 0 -1 170
box -8 -3 64 105
use OR2X1  OR2X1_27
timestamp 1681708930
transform -1 0 1288 0 -1 170
box -8 -3 40 105
use M3_M2  M3_M2_3908
timestamp 1681708930
transform 1 0 1324 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_3860
timestamp 1681708930
transform 1 0 1348 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3898
timestamp 1681708930
transform 1 0 1364 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3899
timestamp 1681708930
transform 1 0 1380 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3909
timestamp 1681708930
transform 1 0 1356 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_3910
timestamp 1681708930
transform 1 0 1372 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_4066
timestamp 1681708930
transform 1 0 1380 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4067
timestamp 1681708930
transform 1 0 1388 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4114
timestamp 1681708930
transform 1 0 1300 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4115
timestamp 1681708930
transform 1 0 1324 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4136
timestamp 1681708930
transform 1 0 1308 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_3925
timestamp 1681708930
transform 1 0 1332 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_4137
timestamp 1681708930
transform 1 0 1332 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_4138
timestamp 1681708930
transform 1 0 1340 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_3945
timestamp 1681708930
transform 1 0 1348 0 1 115
box -3 -3 3 3
use M2_M1  M2_M1_4139
timestamp 1681708930
transform 1 0 1356 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_4151
timestamp 1681708930
transform 1 0 1316 0 1 105
box -2 -2 2 2
use M3_M2  M3_M2_3962
timestamp 1681708930
transform 1 0 1308 0 1 95
box -3 -3 3 3
use INVX2  INVX2_251
timestamp 1681708930
transform 1 0 1288 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_3950
timestamp 1681708930
transform 1 0 1340 0 1 105
box -3 -3 3 3
use NAND3X1  NAND3X1_148
timestamp 1681708930
transform -1 0 1336 0 -1 170
box -8 -3 40 105
use M3_M2  M3_M2_3926
timestamp 1681708930
transform 1 0 1388 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_4152
timestamp 1681708930
transform 1 0 1364 0 1 105
box -2 -2 2 2
use M3_M2  M3_M2_3951
timestamp 1681708930
transform 1 0 1372 0 1 105
box -3 -3 3 3
use NAND3X1  NAND3X1_149
timestamp 1681708930
transform -1 0 1368 0 -1 170
box -8 -3 40 105
use INVX2  INVX2_252
timestamp 1681708930
transform -1 0 1384 0 -1 170
box -9 -3 26 105
use M2_M1  M2_M1_4140
timestamp 1681708930
transform 1 0 1396 0 1 115
box -2 -2 2 2
use FILL  FILL_1508
timestamp 1681708930
transform 1 0 1384 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_3861
timestamp 1681708930
transform 1 0 1420 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3900
timestamp 1681708930
transform 1 0 1428 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_4035
timestamp 1681708930
transform 1 0 1436 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_4068
timestamp 1681708930
transform 1 0 1420 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4069
timestamp 1681708930
transform 1 0 1428 0 1 135
box -2 -2 2 2
use OAI21X1  OAI21X1_121
timestamp 1681708930
transform -1 0 1424 0 -1 170
box -8 -3 34 105
use M2_M1  M2_M1_4116
timestamp 1681708930
transform 1 0 1436 0 1 125
box -2 -2 2 2
use FILL  FILL_1509
timestamp 1681708930
transform 1 0 1424 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_3927
timestamp 1681708930
transform 1 0 1444 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3862
timestamp 1681708930
transform 1 0 1460 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_4036
timestamp 1681708930
transform 1 0 1468 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_4070
timestamp 1681708930
transform 1 0 1460 0 1 135
box -2 -2 2 2
use NOR2X1  NOR2X1_86
timestamp 1681708930
transform 1 0 1432 0 -1 170
box -8 -3 32 105
use M3_M2  M3_M2_3911
timestamp 1681708930
transform 1 0 1468 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_4117
timestamp 1681708930
transform 1 0 1468 0 1 125
box -2 -2 2 2
use FILL  FILL_1510
timestamp 1681708930
transform 1 0 1456 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_4037
timestamp 1681708930
transform 1 0 1492 0 1 145
box -2 -2 2 2
use M3_M2  M3_M2_3901
timestamp 1681708930
transform 1 0 1500 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_4071
timestamp 1681708930
transform 1 0 1484 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_3912
timestamp 1681708930
transform 1 0 1500 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_4072
timestamp 1681708930
transform 1 0 1508 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4073
timestamp 1681708930
transform 1 0 1516 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4118
timestamp 1681708930
transform 1 0 1492 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_3952
timestamp 1681708930
transform 1 0 1492 0 1 105
box -3 -3 3 3
use NOR2X1  NOR2X1_87
timestamp 1681708930
transform 1 0 1464 0 -1 170
box -8 -3 32 105
use M3_M2  M3_M2_3928
timestamp 1681708930
transform 1 0 1516 0 1 125
box -3 -3 3 3
use AOI21X1  AOI21X1_55
timestamp 1681708930
transform -1 0 1520 0 -1 170
box -7 -3 39 105
use FILL  FILL_1511
timestamp 1681708930
transform 1 0 1520 0 -1 170
box -8 -3 16 105
use FILL  FILL_1514
timestamp 1681708930
transform 1 0 1528 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_4119
timestamp 1681708930
transform 1 0 1548 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4120
timestamp 1681708930
transform 1 0 1580 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_3953
timestamp 1681708930
transform 1 0 1548 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_3954
timestamp 1681708930
transform 1 0 1580 0 1 105
box -3 -3 3 3
use FILL  FILL_1515
timestamp 1681708930
transform 1 0 1536 0 -1 170
box -8 -3 16 105
use XNOR2X1  XNOR2X1_55
timestamp 1681708930
transform 1 0 1544 0 -1 170
box -8 -3 64 105
use M2_M1  M2_M1_4074
timestamp 1681708930
transform 1 0 1612 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4075
timestamp 1681708930
transform 1 0 1620 0 1 135
box -2 -2 2 2
use FILL  FILL_1516
timestamp 1681708930
transform 1 0 1600 0 -1 170
box -8 -3 16 105
use FILL  FILL_1517
timestamp 1681708930
transform 1 0 1608 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_3913
timestamp 1681708930
transform 1 0 1628 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_3929
timestamp 1681708930
transform 1 0 1636 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_4121
timestamp 1681708930
transform 1 0 1652 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4141
timestamp 1681708930
transform 1 0 1636 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_3955
timestamp 1681708930
transform 1 0 1636 0 1 105
box -3 -3 3 3
use NAND2X1  NAND2X1_100
timestamp 1681708930
transform 1 0 1616 0 -1 170
box -8 -3 32 105
use M3_M2  M3_M2_3902
timestamp 1681708930
transform 1 0 1684 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_4076
timestamp 1681708930
transform 1 0 1684 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_3930
timestamp 1681708930
transform 1 0 1676 0 1 125
box -3 -3 3 3
use OAI21X1  OAI21X1_122
timestamp 1681708930
transform 1 0 1640 0 -1 170
box -8 -3 34 105
use M2_M1  M2_M1_4142
timestamp 1681708930
transform 1 0 1676 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_4143
timestamp 1681708930
transform 1 0 1684 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_3956
timestamp 1681708930
transform 1 0 1684 0 1 105
box -3 -3 3 3
use FILL  FILL_1518
timestamp 1681708930
transform 1 0 1672 0 -1 170
box -8 -3 16 105
use FILL  FILL_1519
timestamp 1681708930
transform 1 0 1680 0 -1 170
box -8 -3 16 105
use FILL  FILL_1520
timestamp 1681708930
transform 1 0 1688 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_4077
timestamp 1681708930
transform 1 0 1724 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4078
timestamp 1681708930
transform 1 0 1732 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_3931
timestamp 1681708930
transform 1 0 1724 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_4122
timestamp 1681708930
transform 1 0 1732 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4123
timestamp 1681708930
transform 1 0 1748 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4144
timestamp 1681708930
transform 1 0 1708 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_4145
timestamp 1681708930
transform 1 0 1724 0 1 115
box -2 -2 2 2
use FILL  FILL_1530
timestamp 1681708930
transform 1 0 1696 0 -1 170
box -8 -3 16 105
use NAND2X1  NAND2X1_101
timestamp 1681708930
transform -1 0 1728 0 -1 170
box -8 -3 32 105
use M3_M2  M3_M2_3914
timestamp 1681708930
transform 1 0 1764 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_4124
timestamp 1681708930
transform 1 0 1764 0 1 125
box -2 -2 2 2
use OAI21X1  OAI21X1_123
timestamp 1681708930
transform -1 0 1760 0 -1 170
box -8 -3 34 105
use M2_M1  M2_M1_4079
timestamp 1681708930
transform 1 0 1772 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4080
timestamp 1681708930
transform 1 0 1780 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_3932
timestamp 1681708930
transform 1 0 1772 0 1 125
box -3 -3 3 3
use FILL  FILL_1531
timestamp 1681708930
transform 1 0 1760 0 -1 170
box -8 -3 16 105
use FILL  FILL_1532
timestamp 1681708930
transform 1 0 1768 0 -1 170
box -8 -3 16 105
use INVX2  INVX2_257
timestamp 1681708930
transform 1 0 1776 0 -1 170
box -9 -3 26 105
use M2_M1  M2_M1_4081
timestamp 1681708930
transform 1 0 1844 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_3933
timestamp 1681708930
transform 1 0 1820 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_4125
timestamp 1681708930
transform 1 0 1828 0 1 125
box -2 -2 2 2
use XNOR2X1  XNOR2X1_56
timestamp 1681708930
transform 1 0 1792 0 -1 170
box -8 -3 64 105
use FILL  FILL_1533
timestamp 1681708930
transform 1 0 1848 0 -1 170
box -8 -3 16 105
use FILL  FILL_1542
timestamp 1681708930
transform 1 0 1856 0 -1 170
box -8 -3 16 105
use FILL  FILL_1543
timestamp 1681708930
transform 1 0 1864 0 -1 170
box -8 -3 16 105
use FILL  FILL_1544
timestamp 1681708930
transform 1 0 1872 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_4082
timestamp 1681708930
transform 1 0 1900 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_3934
timestamp 1681708930
transform 1 0 1892 0 1 125
box -3 -3 3 3
use FILL  FILL_1545
timestamp 1681708930
transform 1 0 1880 0 -1 170
box -8 -3 16 105
use FILL  FILL_1546
timestamp 1681708930
transform 1 0 1888 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_3935
timestamp 1681708930
transform 1 0 1924 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_4126
timestamp 1681708930
transform 1 0 1932 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4146
timestamp 1681708930
transform 1 0 1956 0 1 115
box -2 -2 2 2
use XNOR2X1  XNOR2X1_60
timestamp 1681708930
transform 1 0 1896 0 -1 170
box -8 -3 64 105
use FILL  FILL_1547
timestamp 1681708930
transform 1 0 1952 0 -1 170
box -8 -3 16 105
use FILL  FILL_1548
timestamp 1681708930
transform 1 0 1960 0 -1 170
box -8 -3 16 105
use FILL  FILL_1549
timestamp 1681708930
transform 1 0 1968 0 -1 170
box -8 -3 16 105
use FILL  FILL_1550
timestamp 1681708930
transform 1 0 1976 0 -1 170
box -8 -3 16 105
use FILL  FILL_1551
timestamp 1681708930
transform 1 0 1984 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_3903
timestamp 1681708930
transform 1 0 2004 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_4083
timestamp 1681708930
transform 1 0 2004 0 1 135
box -2 -2 2 2
use FILL  FILL_1552
timestamp 1681708930
transform 1 0 1992 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_3904
timestamp 1681708930
transform 1 0 2028 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_4084
timestamp 1681708930
transform 1 0 2020 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4085
timestamp 1681708930
transform 1 0 2028 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4127
timestamp 1681708930
transform 1 0 2012 0 1 125
box -2 -2 2 2
use NAND2X1  NAND2X1_106
timestamp 1681708930
transform -1 0 2024 0 -1 170
box -8 -3 32 105
use M3_M2  M3_M2_3915
timestamp 1681708930
transform 1 0 2036 0 1 135
box -3 -3 3 3
use FILL  FILL_1553
timestamp 1681708930
transform 1 0 2024 0 -1 170
box -8 -3 16 105
use FILL  FILL_1554
timestamp 1681708930
transform 1 0 2032 0 -1 170
box -8 -3 16 105
use FILL  FILL_1555
timestamp 1681708930
transform 1 0 2040 0 -1 170
box -8 -3 16 105
use FILL  FILL_1556
timestamp 1681708930
transform 1 0 2048 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_4086
timestamp 1681708930
transform 1 0 2068 0 1 135
box -2 -2 2 2
use FILL  FILL_1557
timestamp 1681708930
transform 1 0 2056 0 -1 170
box -8 -3 16 105
use FILL  FILL_1558
timestamp 1681708930
transform 1 0 2064 0 -1 170
box -8 -3 16 105
use FILL  FILL_1559
timestamp 1681708930
transform 1 0 2072 0 -1 170
box -8 -3 16 105
use FILL  FILL_1560
timestamp 1681708930
transform 1 0 2080 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_4038
timestamp 1681708930
transform 1 0 2100 0 1 145
box -2 -2 2 2
use FILL  FILL_1561
timestamp 1681708930
transform 1 0 2088 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_3916
timestamp 1681708930
transform 1 0 2108 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_4087
timestamp 1681708930
transform 1 0 2116 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_3946
timestamp 1681708930
transform 1 0 2116 0 1 115
box -3 -3 3 3
use M2_M1  M2_M1_4147
timestamp 1681708930
transform 1 0 2124 0 1 115
box -2 -2 2 2
use NOR2X1  NOR2X1_93
timestamp 1681708930
transform 1 0 2096 0 -1 170
box -8 -3 32 105
use FILL  FILL_1562
timestamp 1681708930
transform 1 0 2120 0 -1 170
box -8 -3 16 105
use FILL  FILL_1563
timestamp 1681708930
transform 1 0 2128 0 -1 170
box -8 -3 16 105
use FILL  FILL_1564
timestamp 1681708930
transform 1 0 2136 0 -1 170
box -8 -3 16 105
use FILL  FILL_1565
timestamp 1681708930
transform 1 0 2144 0 -1 170
box -8 -3 16 105
use FILL  FILL_1566
timestamp 1681708930
transform 1 0 2152 0 -1 170
box -8 -3 16 105
use FILL  FILL_1567
timestamp 1681708930
transform 1 0 2160 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_3877
timestamp 1681708930
transform 1 0 2180 0 1 155
box -3 -3 3 3
use FILL  FILL_1568
timestamp 1681708930
transform 1 0 2168 0 -1 170
box -8 -3 16 105
use FILL  FILL_1569
timestamp 1681708930
transform 1 0 2176 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_3936
timestamp 1681708930
transform 1 0 2204 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_4148
timestamp 1681708930
transform 1 0 2204 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_4153
timestamp 1681708930
transform 1 0 2212 0 1 105
box -2 -2 2 2
use NAND3X1  NAND3X1_154
timestamp 1681708930
transform -1 0 2216 0 -1 170
box -8 -3 40 105
use M3_M2  M3_M2_3863
timestamp 1681708930
transform 1 0 2276 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_4039
timestamp 1681708930
transform 1 0 2260 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_4088
timestamp 1681708930
transform 1 0 2236 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4089
timestamp 1681708930
transform 1 0 2244 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_3917
timestamp 1681708930
transform 1 0 2252 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_4128
timestamp 1681708930
transform 1 0 2228 0 1 125
box -2 -2 2 2
use INVX2  INVX2_262
timestamp 1681708930
transform -1 0 2232 0 -1 170
box -9 -3 26 105
use M2_M1  M2_M1_4129
timestamp 1681708930
transform 1 0 2260 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_3937
timestamp 1681708930
transform 1 0 2268 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3918
timestamp 1681708930
transform 1 0 2292 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_4130
timestamp 1681708930
transform 1 0 2276 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4149
timestamp 1681708930
transform 1 0 2268 0 1 115
box -2 -2 2 2
use AOI21X1  AOI21X1_60
timestamp 1681708930
transform 1 0 2232 0 -1 170
box -7 -3 39 105
use M2_M1  M2_M1_4150
timestamp 1681708930
transform 1 0 2292 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_4154
timestamp 1681708930
transform 1 0 2284 0 1 105
box -2 -2 2 2
use M3_M2  M3_M2_3964
timestamp 1681708930
transform 1 0 2292 0 1 75
box -3 -3 3 3
use NAND3X1  NAND3X1_155
timestamp 1681708930
transform 1 0 2264 0 -1 170
box -8 -3 40 105
use FILL  FILL_1570
timestamp 1681708930
transform 1 0 2296 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_3864
timestamp 1681708930
transform 1 0 2316 0 1 165
box -3 -3 3 3
use FILL  FILL_1571
timestamp 1681708930
transform 1 0 2304 0 -1 170
box -8 -3 16 105
use FILL  FILL_1572
timestamp 1681708930
transform 1 0 2312 0 -1 170
box -8 -3 16 105
use FILL  FILL_1573
timestamp 1681708930
transform 1 0 2320 0 -1 170
box -8 -3 16 105
use FILL  FILL_1574
timestamp 1681708930
transform 1 0 2328 0 -1 170
box -8 -3 16 105
use FILL  FILL_1575
timestamp 1681708930
transform 1 0 2336 0 -1 170
box -8 -3 16 105
use FILL  FILL_1576
timestamp 1681708930
transform 1 0 2344 0 -1 170
box -8 -3 16 105
use FILL  FILL_1577
timestamp 1681708930
transform 1 0 2352 0 -1 170
box -8 -3 16 105
use FILL  FILL_1578
timestamp 1681708930
transform 1 0 2360 0 -1 170
box -8 -3 16 105
use FILL  FILL_1579
timestamp 1681708930
transform 1 0 2368 0 -1 170
box -8 -3 16 105
use FILL  FILL_1580
timestamp 1681708930
transform 1 0 2376 0 -1 170
box -8 -3 16 105
use FILL  FILL_1581
timestamp 1681708930
transform 1 0 2384 0 -1 170
box -8 -3 16 105
use FILL  FILL_1582
timestamp 1681708930
transform 1 0 2392 0 -1 170
box -8 -3 16 105
use FILL  FILL_1583
timestamp 1681708930
transform 1 0 2400 0 -1 170
box -8 -3 16 105
use FILL  FILL_1584
timestamp 1681708930
transform 1 0 2408 0 -1 170
box -8 -3 16 105
use FILL  FILL_1585
timestamp 1681708930
transform 1 0 2416 0 -1 170
box -8 -3 16 105
use FILL  FILL_1586
timestamp 1681708930
transform 1 0 2424 0 -1 170
box -8 -3 16 105
use FILL  FILL_1587
timestamp 1681708930
transform 1 0 2432 0 -1 170
box -8 -3 16 105
use FILL  FILL_1588
timestamp 1681708930
transform 1 0 2440 0 -1 170
box -8 -3 16 105
use FILL  FILL_1589
timestamp 1681708930
transform 1 0 2448 0 -1 170
box -8 -3 16 105
use FILL  FILL_1590
timestamp 1681708930
transform 1 0 2456 0 -1 170
box -8 -3 16 105
use FILL  FILL_1591
timestamp 1681708930
transform 1 0 2464 0 -1 170
box -8 -3 16 105
use FILL  FILL_1592
timestamp 1681708930
transform 1 0 2472 0 -1 170
box -8 -3 16 105
use FILL  FILL_1593
timestamp 1681708930
transform 1 0 2480 0 -1 170
box -8 -3 16 105
use FILL  FILL_1594
timestamp 1681708930
transform 1 0 2488 0 -1 170
box -8 -3 16 105
use FILL  FILL_1595
timestamp 1681708930
transform 1 0 2496 0 -1 170
box -8 -3 16 105
use FILL  FILL_1596
timestamp 1681708930
transform 1 0 2504 0 -1 170
box -8 -3 16 105
use FILL  FILL_1597
timestamp 1681708930
transform 1 0 2512 0 -1 170
box -8 -3 16 105
use FILL  FILL_1598
timestamp 1681708930
transform 1 0 2520 0 -1 170
box -8 -3 16 105
use FILL  FILL_1599
timestamp 1681708930
transform 1 0 2528 0 -1 170
box -8 -3 16 105
use FILL  FILL_1600
timestamp 1681708930
transform 1 0 2536 0 -1 170
box -8 -3 16 105
use FILL  FILL_1601
timestamp 1681708930
transform 1 0 2544 0 -1 170
box -8 -3 16 105
use FILL  FILL_1602
timestamp 1681708930
transform 1 0 2552 0 -1 170
box -8 -3 16 105
use FILL  FILL_1603
timestamp 1681708930
transform 1 0 2560 0 -1 170
box -8 -3 16 105
use FILL  FILL_1604
timestamp 1681708930
transform 1 0 2568 0 -1 170
box -8 -3 16 105
use FILL  FILL_1605
timestamp 1681708930
transform 1 0 2576 0 -1 170
box -8 -3 16 105
use FILL  FILL_1606
timestamp 1681708930
transform 1 0 2584 0 -1 170
box -8 -3 16 105
use FILL  FILL_1607
timestamp 1681708930
transform 1 0 2592 0 -1 170
box -8 -3 16 105
use FILL  FILL_1608
timestamp 1681708930
transform 1 0 2600 0 -1 170
box -8 -3 16 105
use FILL  FILL_1609
timestamp 1681708930
transform 1 0 2608 0 -1 170
box -8 -3 16 105
use FILL  FILL_1610
timestamp 1681708930
transform 1 0 2616 0 -1 170
box -8 -3 16 105
use FILL  FILL_1611
timestamp 1681708930
transform 1 0 2624 0 -1 170
box -8 -3 16 105
use FILL  FILL_1612
timestamp 1681708930
transform 1 0 2632 0 -1 170
box -8 -3 16 105
use FILL  FILL_1614
timestamp 1681708930
transform 1 0 2640 0 -1 170
box -8 -3 16 105
use FILL  FILL_1616
timestamp 1681708930
transform 1 0 2648 0 -1 170
box -8 -3 16 105
use FILL  FILL_1618
timestamp 1681708930
transform 1 0 2656 0 -1 170
box -8 -3 16 105
use top_mod_new_VIA0  top_mod_new_VIA0_51
timestamp 1681708930
transform 1 0 2712 0 1 70
box -10 -3 10 3
use top_mod_new_VIA1  top_mod_new_VIA1_4
timestamp 1681708930
transform 1 0 48 0 1 47
box -10 -10 10 10
use top_mod_new_VIA1  top_mod_new_VIA1_5
timestamp 1681708930
transform 1 0 2688 0 1 47
box -10 -10 10 10
use top_mod_new_VIA1  top_mod_new_VIA1_6
timestamp 1681708930
transform 1 0 24 0 1 23
box -10 -10 10 10
use top_mod_new_VIA1  top_mod_new_VIA1_7
timestamp 1681708930
transform 1 0 2712 0 1 23
box -10 -10 10 10
use PadFrame  PadFrame_0
timestamp 1681749783
transform 0 1 1375 -1 0 1300
box -2500 -2500 2500 2500
<< labels >>
rlabel metal3 2 1145 2 1145 4 in_clka
rlabel metal3 2 195 2 195 4 in_clkb
rlabel m3contact 2 1325 2 1325 4 in_restart
rlabel m3contact 2 1005 2 1005 4 in_enable_encode
rlabel metal2 1220 2638 1220 2638 4 in_d_in[6]
rlabel metal2 1148 2638 1148 2638 4 in_d_in[5]
rlabel metal2 1044 2638 1044 2638 4 in_d_in[4]
rlabel metal2 980 2638 980 2638 4 in_d_in[3]
rlabel metal2 852 2638 852 2638 4 in_d_in[2]
rlabel metal2 932 2638 932 2638 4 in_d_in[1]
rlabel metal2 772 2638 772 2638 4 in_d_in[0]
rlabel m3contact 2 2135 2 2135 4 in_key_in[7]
rlabel metal3 2 2335 2 2335 4 in_key_in[6]
rlabel metal3 2 2115 2 2115 4 in_key_in[5]
rlabel m3contact 2 2405 2 2405 4 in_key_in[4]
rlabel metal3 2 2205 2 2205 4 in_key_in[3]
rlabel metal3 2 2185 2 2185 4 in_key_in[2]
rlabel metal3 2 2155 2 2155 4 in_key_in[1]
rlabel metal2 476 2638 476 2638 4 in_key_in[0]
rlabel metal3 2 615 2 615 4 out_data[15]
rlabel m3contact 2 815 2 815 4 out_data[14]
rlabel metal3 2 665 2 665 4 out_data[13]
rlabel metal2 292 1 292 1 4 out_data[12]
rlabel metal2 476 1 476 1 4 out_data[11]
rlabel metal2 676 1 676 1 4 out_data[10]
rlabel metal2 660 1 660 1 4 out_data[9]
rlabel metal2 692 1 692 1 4 out_data[8]
rlabel metal2 644 1 644 1 4 out_data[7]
rlabel m3contact 2 715 2 715 4 out_data[5]
rlabel metal2 460 1 460 1 4 out_data[4]
rlabel m3contact 2 335 2 335 4 out_data[3]
rlabel m3contact 2 535 2 535 4 out_data[2]
rlabel m3contact 2 175 2 175 4 out_data[1]
rlabel metal2 204 1 204 1 4 out_data[0]
rlabel metal1 38 167 38 167 4 gnd
rlabel metal1 14 67 14 67 4 vdd
rlabel metal2 1348 2638 1348 2638 4 in_d_in[7]
rlabel m3contact 2 735 2 735 4 out_data[6]
rlabel pad 1216 -1047 1216 -1047 1 GND!
rlabel pad 3740 860 3740 860 1 Vdd!
rlabel pad 1534 3671 1534 3671 1 GND!
rlabel pad -1001 1460 -1001 1460 1 Vdd!
rlabel pad 3739 1157 3739 1157 1 d_in_7
rlabel pad 3750 1443 3750 1443 1 d_in_6
rlabel pad 3746 1755 3746 1755 1 d_in_5
rlabel pad 3736 2045 3736 2045 1 d_in_4
rlabel pad 3745 2354 3745 2354 1 d_in_3
rlabel pad 3741 2638 3741 2638 1 d_in_1
rlabel pad 2717 3661 2717 3661 1 d_in_2
rlabel pad 2427 3664 2427 3664 1 d_in_0
rlabel pad 2122 3661 2122 3661 1 key_in_0
rlabel pad 1829 3677 1829 3677 1 key_in_4
rlabel pad 1224 3674 1224 3674 1 key_in_6
rlabel pad 933 3666 933 3666 1 key_in_3
rlabel pad 622 3669 622 3669 1 key_in_2
rlabel pad 309 3671 309 3671 1 key_in_1
rlabel pad 20 3673 20 3673 1 key_in_7
rlabel pad -999 2649 -999 2649 1 key_in_5
rlabel pad -995 2354 -995 2354 1 in_restart
rlabel pad -1003 2042 -1003 2042 1 in_clka
rlabel pad -998 1749 -998 1749 1 in_enable_encode
rlabel pad -1015 1137 -1015 1137 1 out_data_14
rlabel pad -1000 841 -1000 841 1 out_data_6
rlabel pad -1006 551 -1006 551 1 out_data_5
rlabel pad -1009 256 -1009 256 1 out_data_13
rlabel pad -1008 -55 -1008 -55 1 out_data_15
rlabel pad 26 -1057 26 -1057 1 out_data_2
rlabel pad 327 -1066 327 -1066 1 out_data_3
rlabel pad 625 -1067 625 -1067 1 out_data_1
rlabel pad 929 -1060 929 -1060 1 in_clkb
rlabel pad 1523 -1066 1523 -1066 1 out_data_0
rlabel pad 1831 -1062 1831 -1062 1 out_data_12
rlabel pad 2123 -1081 2123 -1081 1 out_data_4
rlabel pad 2433 -1080 2433 -1080 1 out_data_11
rlabel pad 2725 -1075 2725 -1075 1 out_data_7
rlabel pad 3743 -51 3743 -51 1 out_data_9
rlabel pad 3739 253 3739 253 1 out_data_10
rlabel pad 3744 555 3744 555 1 out_data_8
<< end >>
