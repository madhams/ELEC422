magic
tech scmos
timestamp 1681708930
<< m2contact >>
rect -2 -2 2 2
<< end >>
